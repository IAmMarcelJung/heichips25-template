module heichips25_tiny_wrapper (clk,
    ena,
    rst_n,
    VPWR,
    VGND,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 inout VPWR;
 inout VGND;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net146;
 wire net147;
 wire net148;
 wire net149;
 wire net150;
 wire net151;
 wire net152;
 wire net153;
 wire net154;
 wire net155;
 wire net156;
 wire net157;
 wire net158;
 wire net159;
 wire net160;
 wire net161;
 wire net162;
 wire net163;
 wire net164;
 wire net165;
 wire net166;
 wire net167;
 wire net168;
 wire net169;
 wire net170;
 wire net171;
 wire net172;
 wire net173;
 wire net174;
 wire net175;
 wire net176;
 wire net177;
 wire net178;
 wire net179;
 wire net180;
 wire net181;
 wire net182;
 wire net183;
 wire net184;
 wire net185;
 wire net186;
 wire net187;
 wire net188;
 wire net189;
 wire net190;
 wire net191;
 wire net192;
 wire net193;
 wire net194;
 wire net195;
 wire net196;
 wire net197;
 wire net198;
 wire net199;
 wire net200;
 wire net201;
 wire net202;
 wire net203;
 wire net204;
 wire net205;
 wire net206;
 wire net207;
 wire net208;
 wire net209;
 wire net210;
 wire net211;
 wire net212;
 wire net213;
 wire net214;
 wire net215;
 wire net216;
 wire net217;
 wire net218;
 wire net219;
 wire net220;
 wire net221;
 wire net222;
 wire net223;
 wire net224;
 wire net225;
 wire net226;
 wire net227;
 wire net228;
 wire net229;
 wire net230;
 wire net231;
 wire net232;
 wire net233;
 wire net234;
 wire net235;
 wire net236;
 wire net237;
 wire net238;
 wire net239;
 wire net240;
 wire net241;
 wire net242;
 wire net243;
 wire net244;
 wire net245;
 wire net246;
 wire net247;
 wire net248;
 wire net249;
 wire net250;
 wire net251;
 wire net252;
 wire net253;
 wire net254;
 wire net255;
 wire net256;
 wire net257;
 wire net258;
 wire net259;
 wire net260;
 wire net261;
 wire net262;
 wire net263;
 wire net264;
 wire net265;
 wire net266;
 wire net267;
 wire net268;
 wire net269;
 wire net270;
 wire net271;
 wire net272;
 wire net273;
 wire net274;
 wire net275;
 wire net276;
 wire net277;
 wire net278;
 wire net279;
 wire net280;
 wire net281;
 wire net282;
 wire net283;
 wire net284;
 wire net285;
 wire net286;
 wire net287;
 wire net288;
 wire net289;
 wire net290;
 wire net291;
 wire net292;
 wire net293;
 wire net294;
 wire net295;
 wire net296;
 wire net297;
 wire net298;
 wire net299;
 wire net300;
 wire net301;
 wire net302;
 wire net303;
 wire net304;
 wire net305;
 wire net306;
 wire net307;
 wire net308;
 wire net309;
 wire net310;
 wire net311;
 wire net312;
 wire net313;
 wire net314;
 wire net315;
 wire net316;
 wire net317;
 wire net318;
 wire net319;
 wire net320;
 wire net321;
 wire net322;
 wire net323;
 wire net324;
 wire net325;
 wire net326;
 wire net327;
 wire net328;
 wire net329;
 wire net330;
 wire net331;
 wire net332;
 wire net333;
 wire net334;
 wire net335;
 wire net336;
 wire net337;
 wire net338;
 wire net339;
 wire net340;
 wire net341;
 wire net342;
 wire net343;
 wire net344;
 wire net345;
 wire net346;
 wire net347;
 wire net348;
 wire net349;
 wire net350;
 wire net351;
 wire net352;
 wire net353;
 wire net354;
 wire net355;
 wire net356;
 wire net357;
 wire net358;
 wire net359;
 wire net360;
 wire net361;
 wire net362;
 wire net363;
 wire net364;
 wire net365;
 wire net366;
 wire net367;
 wire net368;
 wire net369;
 wire net370;
 wire net371;
 wire net372;
 wire clknet_leaf_0_clk;
 wire \falu_i.falutop.alu_data_in[0] ;
 wire \falu_i.falutop.alu_data_in[10] ;
 wire \falu_i.falutop.alu_data_in[11] ;
 wire \falu_i.falutop.alu_data_in[12] ;
 wire \falu_i.falutop.alu_data_in[13] ;
 wire \falu_i.falutop.alu_data_in[14] ;
 wire \falu_i.falutop.alu_data_in[15] ;
 wire \falu_i.falutop.alu_data_in[1] ;
 wire \falu_i.falutop.alu_data_in[2] ;
 wire \falu_i.falutop.alu_data_in[3] ;
 wire \falu_i.falutop.alu_data_in[4] ;
 wire \falu_i.falutop.alu_data_in[5] ;
 wire \falu_i.falutop.alu_data_in[6] ;
 wire \falu_i.falutop.alu_data_in[7] ;
 wire \falu_i.falutop.alu_data_in[8] ;
 wire \falu_i.falutop.alu_data_in[9] ;
 wire \falu_i.falutop.alu_inst.op[0] ;
 wire \falu_i.falutop.alu_inst.op[1] ;
 wire \falu_i.falutop.alu_inst.op[2] ;
 wire \falu_i.falutop.alu_inst.op[3] ;
 wire \falu_i.falutop.data_in[0] ;
 wire \falu_i.falutop.data_in[10] ;
 wire \falu_i.falutop.data_in[11] ;
 wire \falu_i.falutop.data_in[12] ;
 wire \falu_i.falutop.data_in[13] ;
 wire \falu_i.falutop.data_in[14] ;
 wire \falu_i.falutop.data_in[15] ;
 wire \falu_i.falutop.data_in[1] ;
 wire \falu_i.falutop.data_in[2] ;
 wire \falu_i.falutop.data_in[3] ;
 wire \falu_i.falutop.data_in[4] ;
 wire \falu_i.falutop.data_in[5] ;
 wire \falu_i.falutop.data_in[6] ;
 wire \falu_i.falutop.data_in[7] ;
 wire \falu_i.falutop.data_in[8] ;
 wire \falu_i.falutop.data_in[9] ;
 wire \falu_i.falutop.div_inst.a[0] ;
 wire \falu_i.falutop.div_inst.a[1] ;
 wire \falu_i.falutop.div_inst.a[2] ;
 wire \falu_i.falutop.div_inst.a[3] ;
 wire \falu_i.falutop.div_inst.a[4] ;
 wire \falu_i.falutop.div_inst.a[5] ;
 wire \falu_i.falutop.div_inst.a[6] ;
 wire \falu_i.falutop.div_inst.a[7] ;
 wire \falu_i.falutop.div_inst.acc[0] ;
 wire \falu_i.falutop.div_inst.acc[1] ;
 wire \falu_i.falutop.div_inst.acc[2] ;
 wire \falu_i.falutop.div_inst.acc[3] ;
 wire \falu_i.falutop.div_inst.acc[4] ;
 wire \falu_i.falutop.div_inst.acc[5] ;
 wire \falu_i.falutop.div_inst.acc[6] ;
 wire \falu_i.falutop.div_inst.acc[7] ;
 wire \falu_i.falutop.div_inst.acc[8] ;
 wire \falu_i.falutop.div_inst.acc_next[0] ;
 wire \falu_i.falutop.div_inst.b1[0] ;
 wire \falu_i.falutop.div_inst.b1[1] ;
 wire \falu_i.falutop.div_inst.b1[2] ;
 wire \falu_i.falutop.div_inst.b1[3] ;
 wire \falu_i.falutop.div_inst.b1[4] ;
 wire \falu_i.falutop.div_inst.b1[5] ;
 wire \falu_i.falutop.div_inst.b1[6] ;
 wire \falu_i.falutop.div_inst.b1[7] ;
 wire \falu_i.falutop.div_inst.b[0] ;
 wire \falu_i.falutop.div_inst.b[1] ;
 wire \falu_i.falutop.div_inst.b[2] ;
 wire \falu_i.falutop.div_inst.b[3] ;
 wire \falu_i.falutop.div_inst.b[4] ;
 wire \falu_i.falutop.div_inst.b[5] ;
 wire \falu_i.falutop.div_inst.b[6] ;
 wire \falu_i.falutop.div_inst.b[7] ;
 wire \falu_i.falutop.div_inst.busy ;
 wire \falu_i.falutop.div_inst.done ;
 wire \falu_i.falutop.div_inst.i[0] ;
 wire \falu_i.falutop.div_inst.i[1] ;
 wire \falu_i.falutop.div_inst.i[2] ;
 wire \falu_i.falutop.div_inst.quo[0] ;
 wire \falu_i.falutop.div_inst.quo[1] ;
 wire \falu_i.falutop.div_inst.quo[2] ;
 wire \falu_i.falutop.div_inst.quo[3] ;
 wire \falu_i.falutop.div_inst.quo[4] ;
 wire \falu_i.falutop.div_inst.quo[5] ;
 wire \falu_i.falutop.div_inst.quo[6] ;
 wire \falu_i.falutop.div_inst.rem[0] ;
 wire \falu_i.falutop.div_inst.rem[1] ;
 wire \falu_i.falutop.div_inst.rem[2] ;
 wire \falu_i.falutop.div_inst.rem[3] ;
 wire \falu_i.falutop.div_inst.rem[4] ;
 wire \falu_i.falutop.div_inst.rem[5] ;
 wire \falu_i.falutop.div_inst.rem[6] ;
 wire \falu_i.falutop.div_inst.rem[7] ;
 wire \falu_i.falutop.div_inst.start ;
 wire \falu_i.falutop.div_inst.val[0] ;
 wire \falu_i.falutop.div_inst.val[1] ;
 wire \falu_i.falutop.div_inst.val[2] ;
 wire \falu_i.falutop.div_inst.val[3] ;
 wire \falu_i.falutop.div_inst.val[4] ;
 wire \falu_i.falutop.div_inst.val[5] ;
 wire \falu_i.falutop.div_inst.val[6] ;
 wire \falu_i.falutop.div_inst.val[7] ;
 wire \falu_i.falutop.i2c_inst.counter[0] ;
 wire \falu_i.falutop.i2c_inst.counter[1] ;
 wire \falu_i.falutop.i2c_inst.counter[2] ;
 wire \falu_i.falutop.i2c_inst.counter[3] ;
 wire \falu_i.falutop.i2c_inst.counter[4] ;
 wire \falu_i.falutop.i2c_inst.data_in[0] ;
 wire \falu_i.falutop.i2c_inst.data_in[10] ;
 wire \falu_i.falutop.i2c_inst.data_in[11] ;
 wire \falu_i.falutop.i2c_inst.data_in[12] ;
 wire \falu_i.falutop.i2c_inst.data_in[13] ;
 wire \falu_i.falutop.i2c_inst.data_in[14] ;
 wire \falu_i.falutop.i2c_inst.data_in[15] ;
 wire \falu_i.falutop.i2c_inst.data_in[16] ;
 wire \falu_i.falutop.i2c_inst.data_in[17] ;
 wire \falu_i.falutop.i2c_inst.data_in[18] ;
 wire \falu_i.falutop.i2c_inst.data_in[19] ;
 wire \falu_i.falutop.i2c_inst.data_in[1] ;
 wire \falu_i.falutop.i2c_inst.data_in[2] ;
 wire \falu_i.falutop.i2c_inst.data_in[3] ;
 wire \falu_i.falutop.i2c_inst.data_in[4] ;
 wire \falu_i.falutop.i2c_inst.data_in[5] ;
 wire \falu_i.falutop.i2c_inst.data_in[6] ;
 wire \falu_i.falutop.i2c_inst.data_in[7] ;
 wire \falu_i.falutop.i2c_inst.data_in[8] ;
 wire \falu_i.falutop.i2c_inst.data_in[9] ;
 wire \falu_i.falutop.i2c_inst.op[0] ;
 wire \falu_i.falutop.i2c_inst.op[1] ;
 wire \falu_i.falutop.i2c_inst.op[2] ;
 wire \falu_i.falutop.i2c_inst.op[3] ;
 wire \falu_i.falutop.i2c_inst.result[0] ;
 wire \falu_i.falutop.i2c_inst.result[10] ;
 wire \falu_i.falutop.i2c_inst.result[11] ;
 wire \falu_i.falutop.i2c_inst.result[12] ;
 wire \falu_i.falutop.i2c_inst.result[13] ;
 wire \falu_i.falutop.i2c_inst.result[14] ;
 wire \falu_i.falutop.i2c_inst.result[15] ;
 wire \falu_i.falutop.i2c_inst.result[1] ;
 wire \falu_i.falutop.i2c_inst.result[2] ;
 wire \falu_i.falutop.i2c_inst.result[3] ;
 wire \falu_i.falutop.i2c_inst.result[4] ;
 wire \falu_i.falutop.i2c_inst.result[5] ;
 wire \falu_i.falutop.i2c_inst.result[6] ;
 wire \falu_i.falutop.i2c_inst.result[7] ;
 wire \falu_i.falutop.i2c_inst.result[8] ;
 wire \falu_i.falutop.i2c_inst.result[9] ;
 wire \falu_i.falutop.i2c_inst.sda_o ;
 wire \falu_i.falutop.i2c_inst.state[0] ;
 wire \falu_i.falutop.i2c_inst.state[1] ;
 wire \ppwm_i.u_ppwm.data_o ;
 wire \ppwm_i.u_ppwm.global_counter[0] ;
 wire \ppwm_i.u_ppwm.global_counter[10] ;
 wire \ppwm_i.u_ppwm.global_counter[11] ;
 wire \ppwm_i.u_ppwm.global_counter[12] ;
 wire \ppwm_i.u_ppwm.global_counter[13] ;
 wire \ppwm_i.u_ppwm.global_counter[14] ;
 wire \ppwm_i.u_ppwm.global_counter[15] ;
 wire \ppwm_i.u_ppwm.global_counter[16] ;
 wire \ppwm_i.u_ppwm.global_counter[17] ;
 wire \ppwm_i.u_ppwm.global_counter[18] ;
 wire \ppwm_i.u_ppwm.global_counter[19] ;
 wire \ppwm_i.u_ppwm.global_counter[1] ;
 wire \ppwm_i.u_ppwm.global_counter[2] ;
 wire \ppwm_i.u_ppwm.global_counter[3] ;
 wire \ppwm_i.u_ppwm.global_counter[4] ;
 wire \ppwm_i.u_ppwm.global_counter[5] ;
 wire \ppwm_i.u_ppwm.global_counter[6] ;
 wire \ppwm_i.u_ppwm.global_counter[7] ;
 wire \ppwm_i.u_ppwm.global_counter[8] ;
 wire \ppwm_i.u_ppwm.global_counter[9] ;
 wire \ppwm_i.u_ppwm.pc[0] ;
 wire \ppwm_i.u_ppwm.pc[1] ;
 wire \ppwm_i.u_ppwm.pc[2] ;
 wire \ppwm_i.u_ppwm.pc[3] ;
 wire \ppwm_i.u_ppwm.period_start ;
 wire \ppwm_i.u_ppwm.polarity ;
 wire \ppwm_i.u_ppwm.pwm_value[0] ;
 wire \ppwm_i.u_ppwm.pwm_value[1] ;
 wire \ppwm_i.u_ppwm.pwm_value[2] ;
 wire \ppwm_i.u_ppwm.pwm_value[3] ;
 wire \ppwm_i.u_ppwm.pwm_value[4] ;
 wire \ppwm_i.u_ppwm.pwm_value[5] ;
 wire \ppwm_i.u_ppwm.pwm_value[6] ;
 wire \ppwm_i.u_ppwm.pwm_value[7] ;
 wire \ppwm_i.u_ppwm.pwm_value[8] ;
 wire \ppwm_i.u_ppwm.pwm_value[9] ;
 wire \ppwm_i.u_ppwm.u_ex.cmp_flag_q ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[0] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[1] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[2] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[3] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[4] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[5] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[6] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[7] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[8] ;
 wire \ppwm_i.u_ppwm.u_ex.reg_value_q[9] ;
 wire \ppwm_i.u_ppwm.u_ex.state_q[0] ;
 wire \ppwm_i.u_ppwm.u_ex.state_q[1] ;
 wire \ppwm_i.u_ppwm.u_ex.state_q[2] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[0] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[1] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[2] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[3] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[4] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[5] ;
 wire \ppwm_i.u_ppwm.u_mem.bit_count[6] ;
 wire \ppwm_i.u_ppwm.u_mem.clk_prog_sync1 ;
 wire \ppwm_i.u_ppwm.u_mem.clk_prog_sync2 ;
 wire \ppwm_i.u_ppwm.u_mem.clk_prog_sync3 ;
 wire \ppwm_i.u_ppwm.u_mem.data_sync1 ;
 wire \ppwm_i.u_ppwm.u_mem.data_sync2 ;
 wire \ppwm_i.u_ppwm.u_mem.memory[0] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[100] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[101] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[102] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[103] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[104] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[105] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[106] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[107] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[108] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[109] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[10] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[110] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[111] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[11] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[12] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[13] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[14] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[15] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[16] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[17] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[18] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[19] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[1] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[20] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[21] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[22] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[23] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[24] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[25] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[26] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[27] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[28] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[29] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[2] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[30] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[31] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[32] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[33] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[34] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[35] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[36] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[37] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[38] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[39] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[3] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[40] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[41] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[42] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[43] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[44] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[45] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[46] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[47] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[48] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[49] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[4] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[50] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[51] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[52] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[53] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[54] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[55] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[56] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[57] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[58] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[59] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[5] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[60] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[61] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[62] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[63] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[64] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[65] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[66] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[67] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[68] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[69] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[6] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[70] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[71] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[72] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[73] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[74] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[75] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[76] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[77] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[78] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[79] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[7] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[80] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[81] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[82] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[83] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[84] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[85] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[86] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[87] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[88] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[89] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[8] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[90] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[91] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[92] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[93] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[94] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[95] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[96] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[97] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[98] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[99] ;
 wire \ppwm_i.u_ppwm.u_mem.memory[9] ;
 wire \ppwm_i.u_ppwm.u_mem.programming ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[0] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[1] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[2] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[3] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[4] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[5] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[6] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[7] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[8] ;
 wire \ppwm_i.u_ppwm.u_pwm.cmp_value[9] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[0] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[1] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[2] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[3] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[4] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[5] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[6] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[7] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[8] ;
 wire \ppwm_i.u_ppwm.u_pwm.counter[9] ;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net6;
 wire net25;
 wire net26;
 wire net27;
 wire net7;
 wire net28;
 wire net29;
 wire net30;
 wire net563;
 wire net564;
 wire net565;
 wire net566;
 wire net567;
 wire net568;
 wire net569;
 wire net570;
 wire net571;
 wire net572;
 wire net573;
 wire net574;
 wire net575;
 wire net576;
 wire net577;
 wire net578;
 wire net579;
 wire net580;
 wire net581;
 wire net582;
 wire net583;
 wire net584;
 wire net585;
 wire net586;
 wire net587;
 wire net588;
 wire net589;
 wire net590;
 wire net591;
 wire net592;
 wire net593;
 wire net594;
 wire net595;
 wire net596;
 wire net597;
 wire net598;
 wire net599;
 wire net600;
 wire net601;
 wire net602;
 wire net603;
 wire net604;
 wire net605;
 wire net606;
 wire net607;
 wire net608;
 wire net609;
 wire net610;
 wire net611;
 wire net612;
 wire net613;
 wire net614;
 wire net615;
 wire net616;
 wire net617;
 wire net618;
 wire net619;
 wire net620;
 wire net621;
 wire net622;
 wire net623;
 wire net624;
 wire net625;
 wire net626;
 wire net627;
 wire net628;
 wire net629;
 wire net630;
 wire net631;
 wire net632;
 wire net633;
 wire net634;
 wire net635;
 wire net636;
 wire net637;
 wire net638;
 wire net639;
 wire net640;
 wire net641;
 wire net642;
 wire net643;
 wire net644;
 wire net645;
 wire net646;
 wire net647;
 wire net648;
 wire net649;
 wire net650;
 wire net651;
 wire net652;
 wire net653;
 wire net654;
 wire net655;
 wire net656;
 wire net657;
 wire net658;
 wire net659;
 wire net660;
 wire net661;
 wire net662;
 wire net663;
 wire net664;
 wire net665;
 wire net666;
 wire net667;
 wire net668;
 wire net669;
 wire net670;
 wire net671;
 wire net672;
 wire net673;
 wire net674;
 wire net675;
 wire net676;
 wire net677;
 wire net678;
 wire net679;
 wire net680;
 wire net681;
 wire net682;
 wire net683;
 wire net684;
 wire net685;
 wire net686;
 wire net687;
 wire net688;
 wire net689;
 wire net690;
 wire net691;
 wire net692;
 wire net693;
 wire net694;
 wire net695;
 wire net696;
 wire net697;
 wire net698;
 wire net699;
 wire net700;
 wire net701;
 wire net702;
 wire net703;
 wire net704;
 wire net705;
 wire net706;
 wire net707;
 wire net708;
 wire net709;
 wire net710;
 wire net711;
 wire net712;
 wire net713;
 wire net714;
 wire net715;
 wire net716;
 wire net717;
 wire net718;
 wire net719;
 wire net720;
 wire net721;
 wire net722;
 wire net723;
 wire net724;
 wire net725;
 wire net726;
 wire net727;
 wire net728;
 wire net729;
 wire net730;
 wire net731;
 wire net732;
 wire net733;
 wire net734;
 wire net735;
 wire net736;
 wire net737;
 wire net738;
 wire net739;
 wire net740;
 wire net741;
 wire net742;
 wire net743;
 wire net744;
 wire net745;
 wire net746;
 wire net747;
 wire net748;
 wire net749;
 wire net750;
 wire net751;
 wire net752;
 wire net753;
 wire net754;
 wire net755;
 wire net756;
 wire net757;
 wire net758;
 wire net759;
 wire net760;
 wire net761;
 wire net762;
 wire net763;
 wire net764;
 wire net765;
 wire net766;
 wire net767;
 wire net768;
 wire net769;
 wire net770;
 wire net771;
 wire net772;
 wire net773;
 wire net774;
 wire net775;
 wire net776;
 wire net777;
 wire net778;
 wire net779;
 wire net780;
 wire net781;
 wire net782;
 wire net783;
 wire net784;
 wire net785;
 wire net786;
 wire net787;
 wire net788;
 wire net789;
 wire net790;
 wire net791;
 wire net792;
 wire net793;
 wire net794;
 wire net795;
 wire net796;
 wire net797;
 wire net798;
 wire net799;
 wire net800;
 wire net801;
 wire net802;
 wire net803;
 wire net804;
 wire net805;
 wire net806;
 wire net807;
 wire net808;
 wire net809;
 wire net810;
 wire net811;
 wire net812;
 wire net813;
 wire net814;
 wire net815;
 wire net816;
 wire net817;
 wire net818;
 wire net819;
 wire net820;
 wire net821;
 wire net822;
 wire net823;
 wire net824;
 wire net825;
 wire net826;
 wire net827;
 wire net828;
 wire net829;
 wire net830;
 wire net831;
 wire net832;
 wire net833;
 wire net834;
 wire net835;
 wire net836;
 wire net837;
 wire net838;
 wire net839;
 wire net840;
 wire net841;
 wire net842;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net8;
 wire clknet_leaf_1_clk;
 wire clknet_leaf_2_clk;
 wire clknet_leaf_3_clk;
 wire clknet_leaf_4_clk;
 wire clknet_leaf_5_clk;
 wire clknet_leaf_6_clk;
 wire clknet_leaf_7_clk;
 wire clknet_leaf_8_clk;
 wire clknet_leaf_9_clk;
 wire clknet_leaf_10_clk;
 wire clknet_leaf_11_clk;
 wire clknet_leaf_12_clk;
 wire clknet_leaf_13_clk;
 wire clknet_leaf_14_clk;
 wire clknet_leaf_15_clk;
 wire clknet_leaf_16_clk;
 wire clknet_leaf_17_clk;
 wire clknet_leaf_18_clk;
 wire clknet_leaf_19_clk;
 wire clknet_leaf_20_clk;
 wire clknet_leaf_21_clk;
 wire clknet_leaf_22_clk;
 wire clknet_leaf_23_clk;
 wire clknet_leaf_24_clk;
 wire clknet_leaf_25_clk;
 wire clknet_leaf_26_clk;
 wire clknet_leaf_27_clk;
 wire clknet_leaf_28_clk;
 wire clknet_leaf_29_clk;
 wire clknet_leaf_30_clk;
 wire clknet_leaf_31_clk;
 wire clknet_leaf_32_clk;
 wire clknet_leaf_33_clk;
 wire clknet_leaf_34_clk;
 wire clknet_leaf_35_clk;
 wire clknet_leaf_36_clk;
 wire clknet_leaf_37_clk;
 wire clknet_leaf_38_clk;
 wire clknet_leaf_39_clk;
 wire clknet_leaf_40_clk;
 wire clknet_leaf_41_clk;
 wire clknet_leaf_42_clk;
 wire clknet_leaf_43_clk;
 wire clknet_leaf_44_clk;
 wire clknet_0_clk;
 wire clknet_3_0__leaf_clk;
 wire clknet_3_1__leaf_clk;
 wire clknet_3_2__leaf_clk;
 wire clknet_3_3__leaf_clk;
 wire clknet_3_4__leaf_clk;
 wire clknet_3_5__leaf_clk;
 wire clknet_3_6__leaf_clk;
 wire clknet_3_7__leaf_clk;
 wire net373;
 wire net374;
 wire net375;
 wire net376;
 wire net377;
 wire net378;
 wire net379;
 wire net380;
 wire net381;
 wire net382;
 wire net383;
 wire net384;
 wire net385;
 wire net386;
 wire net387;
 wire net388;
 wire net389;
 wire net390;
 wire net391;
 wire net392;
 wire net393;
 wire net394;
 wire net395;
 wire net396;
 wire net397;
 wire net398;
 wire net399;
 wire net400;
 wire net401;
 wire net402;
 wire net403;
 wire net404;
 wire net405;
 wire net406;
 wire net407;
 wire net408;
 wire net409;
 wire net410;
 wire net411;
 wire net412;
 wire net413;
 wire net414;
 wire net415;
 wire net416;
 wire net417;
 wire net418;
 wire net419;
 wire net420;
 wire net421;
 wire net422;
 wire net423;
 wire net424;
 wire net425;
 wire net426;
 wire net427;
 wire net428;
 wire net429;
 wire net430;
 wire net431;
 wire net432;
 wire net433;
 wire net434;
 wire net435;
 wire net436;
 wire net437;
 wire net438;
 wire net439;
 wire net440;
 wire net441;
 wire net442;
 wire net443;
 wire net444;
 wire net445;
 wire net446;
 wire net447;
 wire net448;
 wire net449;
 wire net450;
 wire net451;
 wire net452;
 wire net453;
 wire net454;
 wire net455;
 wire net456;
 wire net457;
 wire net458;
 wire net459;
 wire net460;
 wire net461;
 wire net462;
 wire net463;
 wire net464;
 wire net465;
 wire net466;
 wire net467;
 wire net468;
 wire net469;
 wire net470;
 wire net471;
 wire net472;
 wire net473;
 wire net474;
 wire net475;
 wire net476;
 wire net477;
 wire net478;
 wire net479;
 wire net480;
 wire net481;
 wire net482;
 wire net483;
 wire net484;
 wire net485;
 wire net486;
 wire net487;
 wire net488;
 wire net489;
 wire net490;
 wire net491;
 wire net492;
 wire net493;
 wire net494;
 wire net495;
 wire net496;
 wire net497;
 wire net498;
 wire net499;
 wire net500;
 wire net501;
 wire net502;
 wire net503;
 wire net504;
 wire net505;
 wire net506;
 wire net507;
 wire net508;
 wire net509;
 wire net510;
 wire net511;
 wire net512;
 wire net513;
 wire net514;
 wire net515;
 wire net516;
 wire net517;
 wire net518;
 wire net519;
 wire net520;
 wire net521;
 wire net522;
 wire net523;
 wire net524;
 wire net525;
 wire net526;
 wire net527;
 wire net528;
 wire net529;
 wire net530;
 wire net531;
 wire net532;
 wire net533;
 wire net534;
 wire net535;
 wire net536;
 wire net537;
 wire net538;
 wire net539;
 wire net540;
 wire net541;
 wire net542;
 wire net543;
 wire net544;
 wire net545;
 wire net546;
 wire net547;
 wire net548;
 wire net549;
 wire net550;
 wire net551;
 wire net552;
 wire net553;
 wire net554;
 wire net555;
 wire net556;
 wire net557;
 wire net558;
 wire net559;
 wire net560;
 wire net561;
 wire net562;
 wire net843;
 wire net844;
 wire net845;
 wire net846;
 wire net847;
 wire net848;
 wire net849;
 wire net850;
 wire net851;
 wire net852;
 wire net853;
 wire net854;
 wire net855;
 wire net856;
 wire net857;
 wire net858;
 wire net859;
 wire net860;
 wire net861;
 wire net862;
 wire net863;
 wire net864;
 wire net865;
 wire net866;
 wire net867;
 wire net868;
 wire net869;
 wire net870;
 wire net871;
 wire net872;
 wire net873;
 wire net874;
 wire net875;
 wire net876;
 wire net877;
 wire net878;
 wire net879;
 wire net880;
 wire net881;
 wire net882;
 wire net883;
 wire net884;
 wire net885;
 wire net886;
 wire net887;
 wire net888;
 wire net889;
 wire net890;
 wire net891;
 wire net892;
 wire net893;
 wire net894;
 wire net895;
 wire net896;
 wire net897;
 wire net898;
 wire net899;
 wire net900;
 wire net901;
 wire net902;
 wire net903;
 wire net904;
 wire net905;
 wire net906;
 wire net907;
 wire net908;
 wire net909;
 wire net910;
 wire net911;
 wire net912;
 wire net913;
 wire net914;
 wire net915;
 wire net916;
 wire net917;
 wire net918;
 wire net919;
 wire net920;
 wire net921;
 wire net922;
 wire net923;
 wire net924;
 wire net925;
 wire net926;
 wire net927;
 wire net928;
 wire net929;
 wire net930;
 wire net931;
 wire net932;
 wire net933;
 wire net934;
 wire net935;
 wire net936;
 wire net937;
 wire net938;
 wire net939;
 wire net940;
 wire net941;
 wire net942;
 wire net943;
 wire net944;
 wire net945;
 wire net946;
 wire net947;
 wire net948;
 wire net949;
 wire net950;
 wire net951;
 wire net952;
 wire net953;
 wire net954;
 wire net955;
 wire net956;
 wire net957;
 wire net958;
 wire net959;
 wire net960;
 wire net961;
 wire net962;
 wire net963;
 wire net964;
 wire net965;
 wire net966;
 wire net967;
 wire net968;
 wire net969;
 wire net970;
 wire net971;
 wire net972;
 wire net973;
 wire net974;
 wire net975;
 wire net976;
 wire net977;
 wire net978;
 wire net979;
 wire net980;
 wire net981;
 wire net982;
 wire net983;
 wire net984;
 wire net985;
 wire net986;
 wire net987;
 wire net988;
 wire net989;
 wire net990;
 wire net991;
 wire net992;
 wire net993;
 wire net994;
 wire net995;
 wire net996;
 wire net997;
 wire net998;
 wire net999;
 wire net1000;
 wire net1001;
 wire net1002;
 wire net1003;
 wire net1004;
 wire net1005;
 wire net1006;
 wire net1007;
 wire net1008;
 wire net1009;
 wire net1010;
 wire net1011;
 wire net1012;
 wire net1013;
 wire net1014;
 wire net1015;
 wire net1016;
 wire net1017;
 wire net1018;
 wire net1019;
 wire net1020;
 wire net1021;
 wire net1022;
 wire net1023;
 wire net1024;
 wire net1025;
 wire net1026;
 wire net1027;
 wire net1028;
 wire net1029;
 wire net1030;
 wire net1031;
 wire net1032;
 wire net1033;
 wire net1034;
 wire net1035;
 wire net1036;
 wire net1037;
 wire net1038;
 wire net1039;
 wire net1040;
 wire net1041;
 wire net1042;
 wire net1043;
 wire net1044;
 wire net1045;
 wire net1046;
 wire net1047;
 wire net1048;
 wire net1049;
 wire net1050;
 wire net1051;
 wire net1052;
 wire net1053;
 wire net1054;
 wire net1055;
 wire net1056;
 wire net1057;
 wire net1058;
 wire net1059;
 wire net1060;
 wire net1061;
 wire net1062;
 wire net1063;
 wire net1064;
 wire net1065;
 wire net1066;
 wire net1067;
 wire net1068;
 wire net1069;
 wire net1070;
 wire net1071;
 wire net1072;
 wire net1073;
 wire net1074;
 wire net1075;
 wire net1076;
 wire net1077;
 wire net1078;
 wire net1079;
 wire net1080;
 wire net1081;
 wire net1082;
 wire net1083;
 wire net1084;
 wire net1085;
 wire net1086;
 wire net1087;
 wire net1088;
 wire net1089;
 wire net1090;
 wire net1091;
 wire net1092;
 wire net1093;
 wire net1094;
 wire net1095;
 wire net1096;
 wire net1097;
 wire net1098;
 wire net1099;
 wire net1100;
 wire net1101;
 wire net1102;
 wire net1103;
 wire net1104;
 wire net1105;
 wire net1106;
 wire net1107;
 wire net1108;
 wire net1109;
 wire net1110;
 wire net1111;
 wire net1112;
 wire net1113;
 wire net1114;
 wire net1115;
 wire net1116;
 wire net1117;
 wire net1118;
 wire net1119;
 wire net1120;
 wire net1121;
 wire net1122;
 wire net1123;
 wire net1124;
 wire net1125;
 wire net1126;
 wire net1127;
 wire net1128;
 wire net1129;
 wire net1130;
 wire net1131;
 wire net1132;
 wire net1133;
 wire net1134;
 wire net1135;
 wire net1136;
 wire net1137;
 wire net1138;
 wire net1139;
 wire net1140;
 wire net1141;
 wire net1142;
 wire net1143;
 wire net1144;
 wire net1145;
 wire net1146;
 wire net1147;
 wire net1148;
 wire net1149;
 wire net1150;
 wire net1151;
 wire net1152;
 wire net1153;
 wire net1154;
 wire net1155;
 wire net1156;
 wire net1157;
 wire net1158;
 wire net1159;
 wire net1160;
 wire net1161;
 wire net1162;
 wire net1163;
 wire net1164;
 wire net1165;
 wire net1166;
 wire net1167;
 wire net1168;
 wire net1169;
 wire net1170;
 wire net1171;
 wire net1172;
 wire net1173;
 wire net1174;
 wire net1175;
 wire net1176;
 wire net1177;
 wire net1178;
 wire net1179;
 wire net1180;
 wire net1181;
 wire net1182;
 wire net1183;
 wire net1184;
 wire net1185;
 wire net1186;
 wire net1187;
 wire net1188;
 wire net1189;
 wire net1190;
 wire net1191;
 wire net1192;
 wire net1193;
 wire net1194;
 wire net1195;
 wire net1196;
 wire net1197;

 sg13g2_inv_2 _2792_ (.Y(_2146_),
    .A(net542),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2793_ (.VDD(VPWR),
    .Y(_2147_),
    .A(net432),
    .VSS(VGND));
 sg13g2_inv_1 _2794_ (.VDD(VPWR),
    .Y(_2148_),
    .A(net405),
    .VSS(VGND));
 sg13g2_inv_1 _2795_ (.VDD(VPWR),
    .Y(_2149_),
    .A(net435),
    .VSS(VGND));
 sg13g2_inv_1 _2796_ (.VDD(VPWR),
    .Y(_2150_),
    .A(net411),
    .VSS(VGND));
 sg13g2_inv_1 _2797_ (.VDD(VPWR),
    .Y(_2151_),
    .A(net399),
    .VSS(VGND));
 sg13g2_inv_1 _2798_ (.VDD(VPWR),
    .Y(_2152_),
    .A(net910),
    .VSS(VGND));
 sg13g2_inv_1 _2799_ (.VDD(VPWR),
    .Y(_2153_),
    .A(net409),
    .VSS(VGND));
 sg13g2_inv_2 _2800_ (.Y(_2154_),
    .A(net1006),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2801_ (.VDD(VPWR),
    .Y(_2155_),
    .A(net1051),
    .VSS(VGND));
 sg13g2_inv_1 _2802_ (.VDD(VPWR),
    .Y(_2156_),
    .A(net951),
    .VSS(VGND));
 sg13g2_inv_1 _2803_ (.VDD(VPWR),
    .Y(_2157_),
    .A(net559),
    .VSS(VGND));
 sg13g2_inv_1 _2804_ (.VDD(VPWR),
    .Y(_2158_),
    .A(net461),
    .VSS(VGND));
 sg13g2_inv_1 _2805_ (.VDD(VPWR),
    .Y(_2159_),
    .A(net445),
    .VSS(VGND));
 sg13g2_inv_1 _2806_ (.VDD(VPWR),
    .Y(_2160_),
    .A(net528),
    .VSS(VGND));
 sg13g2_inv_1 _2807_ (.VDD(VPWR),
    .Y(_2161_),
    .A(net914),
    .VSS(VGND));
 sg13g2_inv_2 _2808_ (.Y(_2162_),
    .A(net392),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2809_ (.VDD(VPWR),
    .Y(_2163_),
    .A(net539),
    .VSS(VGND));
 sg13g2_inv_1 _2810_ (.VDD(VPWR),
    .Y(_2164_),
    .A(net500),
    .VSS(VGND));
 sg13g2_inv_1 _2811_ (.VDD(VPWR),
    .Y(_2165_),
    .A(net537),
    .VSS(VGND));
 sg13g2_inv_1 _2812_ (.VDD(VPWR),
    .Y(_2166_),
    .A(net562),
    .VSS(VGND));
 sg13g2_inv_1 _2813_ (.VDD(VPWR),
    .Y(_2167_),
    .A(net532),
    .VSS(VGND));
 sg13g2_inv_1 _2814_ (.VDD(VPWR),
    .Y(_2168_),
    .A(net556),
    .VSS(VGND));
 sg13g2_inv_1 _2815_ (.VDD(VPWR),
    .Y(_2169_),
    .A(net867),
    .VSS(VGND));
 sg13g2_inv_2 _2816_ (.Y(_2170_),
    .A(net390),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2817_ (.VDD(VPWR),
    .Y(_2171_),
    .A(net957),
    .VSS(VGND));
 sg13g2_inv_1 _2818_ (.VDD(VPWR),
    .Y(_2172_),
    .A(net502),
    .VSS(VGND));
 sg13g2_inv_1 _2819_ (.VDD(VPWR),
    .Y(_2173_),
    .A(net518),
    .VSS(VGND));
 sg13g2_inv_1 _2820_ (.VDD(VPWR),
    .Y(_2174_),
    .A(net510),
    .VSS(VGND));
 sg13g2_inv_1 _2821_ (.VDD(VPWR),
    .Y(_2175_),
    .A(net878),
    .VSS(VGND));
 sg13g2_inv_2 _2822_ (.Y(_2176_),
    .A(net417),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2823_ (.VDD(VPWR),
    .Y(_2177_),
    .A(net948),
    .VSS(VGND));
 sg13g2_inv_1 _2824_ (.VDD(VPWR),
    .Y(_2178_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[80] ),
    .VSS(VGND));
 sg13g2_inv_1 _2825_ (.VDD(VPWR),
    .Y(_2179_),
    .A(net545),
    .VSS(VGND));
 sg13g2_inv_1 _2826_ (.VDD(VPWR),
    .Y(_2180_),
    .A(net551),
    .VSS(VGND));
 sg13g2_inv_1 _2827_ (.VDD(VPWR),
    .Y(_2181_),
    .A(net843),
    .VSS(VGND));
 sg13g2_inv_2 _2828_ (.Y(_2182_),
    .A(net383),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2829_ (.VDD(VPWR),
    .Y(_2183_),
    .A(net922),
    .VSS(VGND));
 sg13g2_inv_1 _2830_ (.VDD(VPWR),
    .Y(_2184_),
    .A(net977),
    .VSS(VGND));
 sg13g2_inv_1 _2831_ (.VDD(VPWR),
    .Y(_2185_),
    .A(net415),
    .VSS(VGND));
 sg13g2_inv_1 _2832_ (.VDD(VPWR),
    .Y(_2186_),
    .A(net463),
    .VSS(VGND));
 sg13g2_inv_1 _2833_ (.VDD(VPWR),
    .Y(_2187_),
    .A(net904),
    .VSS(VGND));
 sg13g2_inv_1 _2834_ (.VDD(VPWR),
    .Y(_2188_),
    .A(net889),
    .VSS(VGND));
 sg13g2_inv_1 _2835_ (.VDD(VPWR),
    .Y(_2189_),
    .A(net903),
    .VSS(VGND));
 sg13g2_inv_1 _2836_ (.VDD(VPWR),
    .Y(_2190_),
    .A(net449),
    .VSS(VGND));
 sg13g2_inv_1 _2837_ (.VDD(VPWR),
    .Y(_2191_),
    .A(net491),
    .VSS(VGND));
 sg13g2_inv_1 _2838_ (.VDD(VPWR),
    .Y(_2192_),
    .A(net437),
    .VSS(VGND));
 sg13g2_inv_1 _2839_ (.VDD(VPWR),
    .Y(_2193_),
    .A(net885),
    .VSS(VGND));
 sg13g2_inv_1 _2840_ (.VDD(VPWR),
    .Y(_2194_),
    .A(net866),
    .VSS(VGND));
 sg13g2_inv_1 _2841_ (.VDD(VPWR),
    .Y(_2195_),
    .A(net557),
    .VSS(VGND));
 sg13g2_inv_2 _2842_ (.Y(_2196_),
    .A(net394),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2843_ (.VDD(VPWR),
    .Y(_2197_),
    .A(net469),
    .VSS(VGND));
 sg13g2_inv_1 _2844_ (.VDD(VPWR),
    .Y(_2198_),
    .A(net443),
    .VSS(VGND));
 sg13g2_inv_1 _2845_ (.VDD(VPWR),
    .Y(_2199_),
    .A(net915),
    .VSS(VGND));
 sg13g2_inv_2 _2846_ (.Y(_2200_),
    .A(net407),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2847_ (.VDD(VPWR),
    .Y(_2201_),
    .A(net434),
    .VSS(VGND));
 sg13g2_inv_1 _2848_ (.VDD(VPWR),
    .Y(_2202_),
    .A(net949),
    .VSS(VGND));
 sg13g2_inv_1 _2849_ (.VDD(VPWR),
    .Y(_2203_),
    .A(net530),
    .VSS(VGND));
 sg13g2_inv_1 _2850_ (.VDD(VPWR),
    .Y(_2204_),
    .A(net893),
    .VSS(VGND));
 sg13g2_inv_1 _2851_ (.VDD(VPWR),
    .Y(_2205_),
    .A(net854),
    .VSS(VGND));
 sg13g2_inv_1 _2852_ (.VDD(VPWR),
    .Y(_2206_),
    .A(net969),
    .VSS(VGND));
 sg13g2_inv_1 _2853_ (.VDD(VPWR),
    .Y(_2207_),
    .A(net455),
    .VSS(VGND));
 sg13g2_inv_1 _2854_ (.VDD(VPWR),
    .Y(_2208_),
    .A(net422),
    .VSS(VGND));
 sg13g2_inv_1 _2855_ (.VDD(VPWR),
    .Y(_2209_),
    .A(net424),
    .VSS(VGND));
 sg13g2_inv_1 _2856_ (.VDD(VPWR),
    .Y(_2210_),
    .A(net472),
    .VSS(VGND));
 sg13g2_inv_1 _2857_ (.VDD(VPWR),
    .Y(_2211_),
    .A(net547),
    .VSS(VGND));
 sg13g2_inv_1 _2858_ (.VDD(VPWR),
    .Y(_2212_),
    .A(net534),
    .VSS(VGND));
 sg13g2_inv_1 _2859_ (.VDD(VPWR),
    .Y(_2213_),
    .A(net516),
    .VSS(VGND));
 sg13g2_inv_1 _2860_ (.VDD(VPWR),
    .Y(_2214_),
    .A(net845),
    .VSS(VGND));
 sg13g2_inv_1 _2861_ (.VDD(VPWR),
    .Y(_2215_),
    .A(net959),
    .VSS(VGND));
 sg13g2_inv_1 _2862_ (.VDD(VPWR),
    .Y(_2216_),
    .A(net508),
    .VSS(VGND));
 sg13g2_inv_1 _2863_ (.VDD(VPWR),
    .Y(_2217_),
    .A(net950),
    .VSS(VGND));
 sg13g2_inv_1 _2864_ (.VDD(VPWR),
    .Y(_2218_),
    .A(net402),
    .VSS(VGND));
 sg13g2_inv_1 _2865_ (.VDD(VPWR),
    .Y(_2219_),
    .A(net477),
    .VSS(VGND));
 sg13g2_inv_1 _2866_ (.VDD(VPWR),
    .Y(_2220_),
    .A(net965),
    .VSS(VGND));
 sg13g2_inv_1 _2867_ (.VDD(VPWR),
    .Y(_2221_),
    .A(net875),
    .VSS(VGND));
 sg13g2_inv_1 _2868_ (.VDD(VPWR),
    .Y(_2222_),
    .A(net898),
    .VSS(VGND));
 sg13g2_inv_1 _2869_ (.VDD(VPWR),
    .Y(_2223_),
    .A(net447),
    .VSS(VGND));
 sg13g2_inv_1 _2870_ (.VDD(VPWR),
    .Y(_2224_),
    .A(net496),
    .VSS(VGND));
 sg13g2_inv_2 _2871_ (.Y(_2225_),
    .A(net928),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2872_ (.VDD(VPWR),
    .Y(_2226_),
    .A(net896),
    .VSS(VGND));
 sg13g2_inv_1 _2873_ (.VDD(VPWR),
    .Y(_2227_),
    .A(net888),
    .VSS(VGND));
 sg13g2_inv_1 _2874_ (.VDD(VPWR),
    .Y(_2228_),
    .A(net504),
    .VSS(VGND));
 sg13g2_inv_1 _2875_ (.VDD(VPWR),
    .Y(_2229_),
    .A(net441),
    .VSS(VGND));
 sg13g2_inv_1 _2876_ (.VDD(VPWR),
    .Y(_2230_),
    .A(net451),
    .VSS(VGND));
 sg13g2_inv_1 _2877_ (.VDD(VPWR),
    .Y(_2231_),
    .A(net483),
    .VSS(VGND));
 sg13g2_inv_1 _2878_ (.VDD(VPWR),
    .Y(_2232_),
    .A(net560),
    .VSS(VGND));
 sg13g2_inv_1 _2879_ (.VDD(VPWR),
    .Y(_2233_),
    .A(net852),
    .VSS(VGND));
 sg13g2_inv_1 _2880_ (.VDD(VPWR),
    .Y(_2234_),
    .A(net523),
    .VSS(VGND));
 sg13g2_inv_2 _2881_ (.Y(_2235_),
    .A(net1160),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2882_ (.Y(_2236_),
    .A(net1169),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2883_ (.Y(_2237_),
    .A(net1172),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2884_ (.Y(_2238_),
    .A(net1174),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2885_ (.Y(_2239_),
    .A(net1183),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2886_ (.Y(_2240_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2887_ (.A(net1143),
    .Y(_2241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2888_ (.A(net1144),
    .Y(_2242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2889_ (.Y(_2243_),
    .A(\ppwm_i.u_ppwm.pwm_value[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2890_ (.A(net1176),
    .Y(_2244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2891_ (.Y(_2245_),
    .A(net1190),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2892_ (.A(net1187),
    .Y(_2246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2893_ (.A(net1188),
    .Y(_2247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2894_ (.A(\ppwm_i.u_ppwm.pwm_value[4] ),
    .Y(_2248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2895_ (.A(net1166),
    .Y(_2249_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2896_ (.Y(_2250_),
    .A(\ppwm_i.u_ppwm.pwm_value[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2897_ (.Y(_2251_),
    .A(net1165),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2898_ (.VDD(VPWR),
    .Y(_2252_),
    .A(net376),
    .VSS(VGND));
 sg13g2_inv_2 _2899_ (.Y(_2253_),
    .A(net1162),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2900_ (.A(net786),
    .Y(_2254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2901_ (.Y(_2255_),
    .A(net419),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2902_ (.VDD(VPWR),
    .Y(_2256_),
    .A(net789),
    .VSS(VGND));
 sg13g2_inv_1 _2903_ (.VDD(VPWR),
    .Y(_2257_),
    .A(net793),
    .VSS(VGND));
 sg13g2_inv_2 _2904_ (.Y(_2258_),
    .A(net1031),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2905_ (.Y(_2259_),
    .A(net1076),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2906_ (.VDD(VPWR),
    .Y(_2260_),
    .A(\ppwm_i.u_ppwm.global_counter[17] ),
    .VSS(VGND));
 sg13g2_inv_1 _2907_ (.VDD(VPWR),
    .Y(_2261_),
    .A(\ppwm_i.u_ppwm.global_counter[16] ),
    .VSS(VGND));
 sg13g2_inv_2 _2908_ (.Y(_2262_),
    .A(net1180),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2909_ (.VDD(VPWR),
    .Y(_2263_),
    .A(\ppwm_i.u_ppwm.global_counter[14] ),
    .VSS(VGND));
 sg13g2_inv_1 _2910_ (.VDD(VPWR),
    .Y(_2264_),
    .A(\ppwm_i.u_ppwm.global_counter[13] ),
    .VSS(VGND));
 sg13g2_inv_1 _2911_ (.VDD(VPWR),
    .Y(_2265_),
    .A(\ppwm_i.u_ppwm.global_counter[12] ),
    .VSS(VGND));
 sg13g2_inv_2 _2912_ (.Y(_2266_),
    .A(\ppwm_i.u_ppwm.global_counter[11] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2913_ (.Y(_2267_),
    .A(net553),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2914_ (.Y(_2268_),
    .A(net1092),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2915_ (.Y(_2269_),
    .A(net1184),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2916_ (.Y(_2270_),
    .A(net1107),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2917_ (.Y(_2271_),
    .A(net1189),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2918_ (.Y(_2272_),
    .A(net1003),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2919_ (.Y(_2273_),
    .A(net1024),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2920_ (.VDD(VPWR),
    .Y(_2274_),
    .A(net1094),
    .VSS(VGND));
 sg13g2_inv_1 _2921_ (.VDD(VPWR),
    .Y(_2275_),
    .A(net1066),
    .VSS(VGND));
 sg13g2_inv_1 _2922_ (.VDD(VPWR),
    .Y(_2276_),
    .A(net1060),
    .VSS(VGND));
 sg13g2_inv_1 _2923_ (.VDD(VPWR),
    .Y(_2277_),
    .A(net1090),
    .VSS(VGND));
 sg13g2_inv_1 _2924_ (.VDD(VPWR),
    .Y(_2278_),
    .A(net863),
    .VSS(VGND));
 sg13g2_inv_1 _2925_ (.VDD(VPWR),
    .Y(_2279_),
    .A(net535),
    .VSS(VGND));
 sg13g2_inv_1 _2926_ (.VDD(VPWR),
    .Y(_2280_),
    .A(net924),
    .VSS(VGND));
 sg13g2_inv_2 _2927_ (.Y(_2281_),
    .A(net430),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2928_ (.VDD(VPWR),
    .Y(_2282_),
    .A(net492),
    .VSS(VGND));
 sg13g2_inv_1 _2929_ (.VDD(VPWR),
    .Y(_2283_),
    .A(net426),
    .VSS(VGND));
 sg13g2_inv_1 _2930_ (.VDD(VPWR),
    .Y(_2284_),
    .A(net470),
    .VSS(VGND));
 sg13g2_inv_1 _2931_ (.VDD(VPWR),
    .Y(_2285_),
    .A(net457),
    .VSS(VGND));
 sg13g2_inv_1 _2932_ (.VDD(VPWR),
    .Y(_2286_),
    .A(net520),
    .VSS(VGND));
 sg13g2_inv_1 _2933_ (.VDD(VPWR),
    .Y(_2287_),
    .A(net506),
    .VSS(VGND));
 sg13g2_inv_1 _2934_ (.VDD(VPWR),
    .Y(_2288_),
    .A(net381),
    .VSS(VGND));
 sg13g2_inv_2 _2935_ (.Y(_2289_),
    .A(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2936_ (.VDD(VPWR),
    .Y(_2290_),
    .A(net485),
    .VSS(VGND));
 sg13g2_inv_2 _2937_ (.Y(_2291_),
    .A(net420),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2938_ (.Y(_2292_),
    .A(net428),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2939_ (.Y(_2293_),
    .A(net467),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2940_ (.Y(_2294_),
    .A(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2941_ (.Y(_2295_),
    .A(net740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2942_ (.A(net721),
    .Y(_2296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2943_ (.A(net716),
    .Y(_2297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2944_ (.VDD(VPWR),
    .Y(_2298_),
    .A(net877),
    .VSS(VGND));
 sg13g2_inv_2 _2945_ (.Y(_2299_),
    .A(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2946_ (.Y(_2300_),
    .A(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _2947_ (.A(net769),
    .Y(_2301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2948_ (.VDD(VPWR),
    .Y(_2302_),
    .A(\falu_i.falutop.alu_data_in[7] ),
    .VSS(VGND));
 sg13g2_inv_1 _2949_ (.VDD(VPWR),
    .Y(_2303_),
    .A(net754),
    .VSS(VGND));
 sg13g2_inv_4 _2950_ (.A(net766),
    .Y(_2304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _2951_ (.Y(_2305_),
    .A(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2952_ (.A(net791),
    .B(net793),
    .X(_2306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2953_ (.Y(_2307_),
    .A(net791),
    .B(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2954_ (.B(net788),
    .C(net700),
    .A(net786),
    .Y(_2308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2955_ (.A(net792),
    .B(net793),
    .Y(_2309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _2956_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2310_),
    .B(net794),
    .A(net792));
 sg13g2_nor2b_2 _2957_ (.A(net794),
    .B_N(net792),
    .Y(_2311_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _2958_ (.A(net792),
    .B_N(net794),
    .Y(_2312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _2959_ (.Y(_2313_),
    .B(net794),
    .A_N(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2960_ (.Y(_2314_),
    .B1(net690),
    .B2(_2170_),
    .A2(net702),
    .A1(_2160_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2961_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2165_),
    .C1(net708),
    .B1(net694),
    .A1(_2174_),
    .Y(_2315_),
    .A2(net697));
 sg13g2_and2_1 _2962_ (.A(_2314_),
    .B(_2315_),
    .X(_2316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _2963_ (.A(\ppwm_i.u_ppwm.u_mem.memory[57] ),
    .B(_2310_),
    .Y(_2317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2964_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2190_),
    .A2(net691),
    .Y(_2318_),
    .B1(net789));
 sg13g2_a22oi_1 _2965_ (.Y(_2319_),
    .B1(net695),
    .B2(_2185_),
    .A2(net703),
    .A1(_2180_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _2966_ (.Y(_2320_),
    .A(_2318_),
    .B(_2319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2967_ (.B1(net787),
    .VDD(VPWR),
    .Y(_2321_),
    .VSS(VGND),
    .A1(_2317_),
    .A2(_2320_));
 sg13g2_a22oi_1 _2968_ (.Y(_2322_),
    .B1(net693),
    .B2(_2224_),
    .A2(net701),
    .A1(_2219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2969_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2229_),
    .C1(net789),
    .B1(net689),
    .A1(_2234_),
    .Y(_2323_),
    .A2(net698));
 sg13g2_o21ai_1 _2970_ (.B1(net790),
    .VDD(VPWR),
    .Y(_2324_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[29] ),
    .A2(_2310_));
 sg13g2_a22oi_1 _2971_ (.Y(_2325_),
    .B1(net693),
    .B2(_2205_),
    .A2(net701),
    .A1(_2200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _2972_ (.B1(_2325_),
    .VDD(VPWR),
    .Y(_2326_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[36] ),
    .A2(_2313_));
 sg13g2_a21oi_1 _2973_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2322_),
    .A2(_2323_),
    .Y(_2327_),
    .B1(net787));
 sg13g2_o21ai_1 _2974_ (.B1(_2327_),
    .VDD(VPWR),
    .Y(_2328_),
    .VSS(VGND),
    .A1(_2324_),
    .A2(_2326_));
 sg13g2_o21ai_1 _2975_ (.B1(_2328_),
    .VDD(VPWR),
    .Y(_2329_),
    .VSS(VGND),
    .A1(_2316_),
    .A2(_2321_));
 sg13g2_inv_1 _2976_ (.VDD(VPWR),
    .Y(_2330_),
    .A(_2329_),
    .VSS(VGND));
 sg13g2_nand2_1 _2977_ (.Y(_2331_),
    .A(_2171_),
    .B(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2166_),
    .A2(net694),
    .Y(_2332_),
    .B1(net709));
 sg13g2_a22oi_1 _2979_ (.Y(_2333_),
    .B1(net697),
    .B2(_2175_),
    .A2(net702),
    .A1(_2161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2980_ (.B(_2332_),
    .C(_2333_),
    .A(_2331_),
    .Y(_2334_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2981_ (.Y(_2335_),
    .B1(net695),
    .B2(_2186_),
    .A2(net703),
    .A1(_2181_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2982_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2191_),
    .C1(net789),
    .B1(net691),
    .A1(_2196_),
    .Y(_2336_),
    .A2(net698));
 sg13g2_a21oi_1 _2983_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2335_),
    .A2(_2336_),
    .Y(_2337_),
    .B1(_2254_));
 sg13g2_nor2_1 _2984_ (.A(\ppwm_i.u_ppwm.u_mem.memory[0] ),
    .B(_2310_),
    .Y(_2338_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2985_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2230_),
    .A2(net688),
    .Y(_2339_),
    .B1(net788));
 sg13g2_a221oi_1 _2986_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2225_),
    .C1(_2338_),
    .B1(net693),
    .A1(_2220_),
    .Y(_2340_),
    .A2(net704));
 sg13g2_a22oi_1 _2987_ (.Y(_2341_),
    .B1(net692),
    .B2(_2206_),
    .A2(net696),
    .A1(_2215_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2988_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2210_),
    .C1(net708),
    .B1(net688),
    .A1(_2201_),
    .Y(_2342_),
    .A2(net701));
 sg13g2_a221oi_1 _2989_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2342_),
    .C1(net787),
    .B1(_2341_),
    .A1(_2339_),
    .Y(_2343_),
    .A2(_2340_));
 sg13g2_a21o_2 _2990_ (.A2(_2337_),
    .A1(_2334_),
    .B1(_2343_),
    .X(_2344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _2991_ (.A(_2329_),
    .B(_2344_),
    .X(_2345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _2992_ (.VDD(VPWR),
    .Y(_2346_),
    .A(_2345_),
    .VSS(VGND));
 sg13g2_nand2_1 _2993_ (.Y(_2347_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[72] ),
    .B(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _2994_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[65] ),
    .A2(net691),
    .Y(_2348_),
    .B1(net789));
 sg13g2_a22oi_1 _2995_ (.Y(_2349_),
    .B1(net698),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[58] ),
    .A2(net703),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[79] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _2996_ (.B(_2348_),
    .C(_2349_),
    .A(_2347_),
    .Y(_2350_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _2997_ (.Y(_2351_),
    .B1(net690),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[93] ),
    .A2(net702),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[107] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _2998_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .C1(net709),
    .B1(net694),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .Y(_2352_),
    .A2(net698));
 sg13g2_a21oi_1 _2999_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2351_),
    .A2(_2352_),
    .Y(_2353_),
    .B1(_2254_));
 sg13g2_and2_1 _3000_ (.A(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .B(net693),
    .X(_2354_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3001_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .A2(net689),
    .Y(_2355_),
    .B1(net789));
 sg13g2_a221oi_1 _3002_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[2] ),
    .C1(_2354_),
    .B1(net699),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .Y(_2356_),
    .A2(net701));
 sg13g2_a22oi_1 _3003_ (.Y(_2357_),
    .B1(net689),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[37] ),
    .A2(net696),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3004_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[44] ),
    .C1(net708),
    .B1(net692),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .Y(_2358_),
    .A2(net701));
 sg13g2_a221oi_1 _3005_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2358_),
    .C1(net787),
    .B1(_2357_),
    .A1(_2355_),
    .Y(_2359_),
    .A2(_2356_));
 sg13g2_a21o_2 _3006_ (.A2(_2353_),
    .A1(_2350_),
    .B1(_2359_),
    .X(_2360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3007_ (.A(_2346_),
    .B(_2360_),
    .Y(_2361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3008_ (.Y(_2362_),
    .B1(net697),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .A2(net702),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[111] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3009_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .C1(net709),
    .B1(net690),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[104] ),
    .Y(_2363_),
    .A2(net694));
 sg13g2_nand2_1 _3010_ (.Y(_2364_),
    .A(\ppwm_i.u_ppwm.u_mem.memory[83] ),
    .B(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3011_ (.A2(net691),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .B1(net789),
    .X(_2365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3012_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[76] ),
    .C1(_2365_),
    .B1(net694),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[62] ),
    .Y(_2366_),
    .A2(net697));
 sg13g2_a22oi_1 _3013_ (.Y(_2367_),
    .B1(_2364_),
    .B2(_2366_),
    .A2(_2363_),
    .A1(_2362_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3014_ (.Y(_2368_),
    .B1(net688),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .A2(net700),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3015_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .C1(net788),
    .B1(net692),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[6] ),
    .Y(_2369_),
    .A2(net696));
 sg13g2_and2_1 _3016_ (.A(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .B(net688),
    .X(_2370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3017_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[48] ),
    .A2(net692),
    .Y(_2371_),
    .B1(net708));
 sg13g2_a221oi_1 _3018_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .C1(_2370_),
    .B1(net696),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[55] ),
    .Y(_2372_),
    .A2(net700));
 sg13g2_a221oi_1 _3019_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2372_),
    .C1(net786),
    .B1(_2371_),
    .A1(_2368_),
    .Y(_2373_),
    .A2(_2369_));
 sg13g2_a21o_1 _3020_ (.A2(_2367_),
    .A1(net786),
    .B1(_2373_),
    .X(_2374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_2 _3021_ (.Y(_2375_),
    .A(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3022_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2167_),
    .A2(net690),
    .Y(_2376_),
    .B1(net709));
 sg13g2_nor3_1 _3023_ (.A(\ppwm_i.u_ppwm.u_mem.memory[89] ),
    .B(net792),
    .C(net794),
    .Y(_2377_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3024_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2162_),
    .C1(_2377_),
    .B1(net695),
    .A1(_2157_),
    .Y(_2378_),
    .A2(net702));
 sg13g2_a22oi_1 _3025_ (.Y(_2379_),
    .B1(net694),
    .B2(_2182_),
    .A2(net703),
    .A1(_2176_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3026_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2187_),
    .C1(net789),
    .B1(net690),
    .A1(_2192_),
    .Y(_2380_),
    .A2(net697));
 sg13g2_a221oi_1 _3027_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2380_),
    .C1(_2254_),
    .B1(_2379_),
    .A1(_2376_),
    .Y(_2381_),
    .A2(_2378_));
 sg13g2_nor3_1 _3028_ (.A(\ppwm_i.u_ppwm.u_mem.memory[33] ),
    .B(net791),
    .C(net793),
    .Y(_2382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3029_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2207_),
    .A2(net688),
    .Y(_2383_),
    .B1(net708));
 sg13g2_a221oi_1 _3030_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2202_),
    .C1(_2382_),
    .B1(net692),
    .A1(_2197_),
    .Y(_2384_),
    .A2(net700));
 sg13g2_a21oi_1 _3031_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2221_),
    .A2(net692),
    .Y(_2385_),
    .B1(net788));
 sg13g2_nor3_1 _3032_ (.A(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .B(net791),
    .C(net793),
    .Y(_2386_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3033_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2226_),
    .C1(_2386_),
    .B1(net688),
    .A1(_2216_),
    .Y(_2387_),
    .A2(net700));
 sg13g2_a221oi_1 _3034_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2387_),
    .C1(net786),
    .B1(_2385_),
    .A1(_2383_),
    .Y(_2388_),
    .A2(_2384_));
 sg13g2_nor2_1 _3035_ (.A(_2381_),
    .B(_2388_),
    .Y(_2389_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3036_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_2390_),
    .B(net612),
    .A(net603));
 sg13g2_nand2b_1 _3037_ (.Y(_2391_),
    .B(net702),
    .A_N(\ppwm_i.u_ppwm.u_mem.memory[108] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3038_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2164_),
    .A2(net694),
    .Y(_2392_),
    .B1(net709));
 sg13g2_a22oi_1 _3039_ (.Y(_2393_),
    .B1(net690),
    .B2(_2169_),
    .A2(net697),
    .A1(_2173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3040_ (.B(_2392_),
    .C(_2393_),
    .A(_2391_),
    .Y(_2394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3041_ (.Y(_2395_),
    .B1(net691),
    .B2(_2189_),
    .A2(net694),
    .A1(_2184_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3042_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2194_),
    .C1(net790),
    .B1(net697),
    .A1(_2178_),
    .Y(_2396_),
    .A2(net703));
 sg13g2_a21oi_1 _3043_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2395_),
    .A2(_2396_),
    .Y(_2397_),
    .B1(_2254_));
 sg13g2_a21oi_1 _3044_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2199_),
    .A2(net704),
    .Y(_2398_),
    .B1(net708));
 sg13g2_nor2_1 _3045_ (.A(\ppwm_i.u_ppwm.u_mem.memory[38] ),
    .B(_2313_),
    .Y(_2399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3046_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2204_),
    .C1(_2399_),
    .B1(net693),
    .A1(_2213_),
    .Y(_2400_),
    .A2(net699));
 sg13g2_a22oi_1 _3047_ (.Y(_2401_),
    .B1(net693),
    .B2(_2223_),
    .A2(net701),
    .A1(_2218_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3048_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2228_),
    .C1(net790),
    .B1(net689),
    .A1(_2233_),
    .Y(_2402_),
    .A2(net696));
 sg13g2_a221oi_1 _3049_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2402_),
    .C1(net787),
    .B1(_2401_),
    .A1(_2398_),
    .Y(_2403_),
    .A2(_2400_));
 sg13g2_a21oi_2 _3050_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2403_),
    .Y(_2404_),
    .A2(_2397_),
    .A1(_2394_));
 sg13g2_nor3_1 _3051_ (.A(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .B(net792),
    .C(net794),
    .Y(_2405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3052_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2168_),
    .A2(net690),
    .Y(_2406_),
    .B1(net709));
 sg13g2_a221oi_1 _3053_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2163_),
    .C1(_2405_),
    .B1(net695),
    .A1(_2158_),
    .Y(_2407_),
    .A2(net702));
 sg13g2_a22oi_1 _3054_ (.Y(_2408_),
    .B1(net691),
    .B2(_2188_),
    .A2(net697),
    .A1(_2193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3055_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2183_),
    .C1(net790),
    .B1(net695),
    .A1(_2177_),
    .Y(_2409_),
    .A2(net703));
 sg13g2_a22oi_1 _3056_ (.Y(_2410_),
    .B1(_2408_),
    .B2(_2409_),
    .A2(_2407_),
    .A1(_2406_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3057_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2208_),
    .A2(net688),
    .Y(_2411_),
    .B1(net708));
 sg13g2_nand2_1 _3058_ (.Y(_2412_),
    .A(_2203_),
    .B(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3059_ (.Y(_2413_),
    .B1(net696),
    .B2(_2212_),
    .A2(net700),
    .A1(_2198_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3060_ (.B(_2412_),
    .C(_2413_),
    .A(_2411_),
    .Y(_2414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3061_ (.Y(_2415_),
    .B1(net692),
    .B2(_2222_),
    .A2(net700),
    .A1(_2217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3062_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2227_),
    .C1(net790),
    .B1(net688),
    .A1(_2232_),
    .Y(_2416_),
    .A2(net696));
 sg13g2_a21oi_1 _3063_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2415_),
    .A2(_2416_),
    .Y(_2417_),
    .B1(net786));
 sg13g2_a22oi_1 _3064_ (.Y(_2418_),
    .B1(_2414_),
    .B2(_2417_),
    .A2(_2410_),
    .A1(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 _3065_ (.A(net608),
    .Y(_2419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3066_ (.A(net585),
    .B(net608),
    .Y(_2420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3067_ (.B(net598),
    .C(_2420_),
    .A(_2361_),
    .Y(_2421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3068_ (.Y(_2422_),
    .A(net419),
    .B(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3069_ (.A(_2422_),
    .B_N(_2421_),
    .Y(_2423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3070_ (.Y(_2424_),
    .B(_2423_),
    .A_N(_2308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3071_ (.Y(_2425_),
    .B(net980),
    .A_N(\ppwm_i.u_ppwm.period_start ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3072_ (.B(_2424_),
    .C(net981),
    .A(net821),
    .Y(_0000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3073_ (.B(net821),
    .C(net385),
    .Y(_2426_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\ppwm_i.u_ppwm.period_start ));
 sg13g2_o21ai_1 _3074_ (.B1(net386),
    .VDD(VPWR),
    .Y(_0001_),
    .VSS(VGND),
    .A1(_2421_),
    .A2(_2422_));
 sg13g2_nand2_1 _3075_ (.Y(_2427_),
    .A(_2308_),
    .B(_2423_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3076_ (.A(net980),
    .B(net385),
    .Y(_2428_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3077_ (.Y(_2429_),
    .A(net1039),
    .B(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3078_ (.B1(_2427_),
    .VDD(VPWR),
    .Y(_0002_),
    .VSS(VGND),
    .A1(_2428_),
    .A2(_2429_));
 sg13g2_nor2_2 _3079_ (.A(net985),
    .B(net1013),
    .Y(_2430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3080_ (.Y(_2431_),
    .A(net1016),
    .B(_2430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3081_ (.A(\falu_i.falutop.i2c_inst.counter[1] ),
    .B(\falu_i.falutop.i2c_inst.counter[0] ),
    .X(_2432_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3082_ (.A(net1001),
    .B_N(\falu_i.falutop.i2c_inst.state[0] ),
    .Y(_2433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3083_ (.Y(_2434_),
    .A(_2432_),
    .B(_2433_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3084_ (.A(_2431_),
    .B(_2434_),
    .Y(_2435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3085_ (.B1(net820),
    .VDD(VPWR),
    .Y(_2436_),
    .VSS(VGND),
    .A1(net1069),
    .A2(_2435_));
 sg13g2_a21oi_1 _3086_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_2435_),
    .Y(_0003_),
    .B1(_2436_));
 sg13g2_nand2b_2 _3087_ (.Y(_2437_),
    .B(_2430_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net1150));
 sg13g2_nor2_2 _3088_ (.A(\falu_i.falutop.i2c_inst.counter[1] ),
    .B(net1045),
    .Y(_2438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3089_ (.Y(_2439_),
    .A(_2433_),
    .B(_2438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3090_ (.A(net1097),
    .B(\falu_i.falutop.i2c_inst.counter[1] ),
    .C(net1045),
    .Y(_2440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3091_ (.A(net985),
    .B_N(_2440_),
    .Y(_2441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3092_ (.Y(_2442_),
    .B(_2438_),
    .A_N(_2437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3093_ (.A(net1014),
    .B(_2439_),
    .Y(_2443_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3094_ (.B1(net816),
    .VDD(VPWR),
    .Y(_2444_),
    .VSS(VGND),
    .A1(net848),
    .A2(_2443_));
 sg13g2_a21oi_1 _3095_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_2443_),
    .Y(_0004_),
    .B1(_2444_));
 sg13g2_nor2b_2 _3096_ (.A(\falu_i.falutop.i2c_inst.counter[1] ),
    .B_N(\falu_i.falutop.i2c_inst.counter[0] ),
    .Y(_2445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3097_ (.Y(_2446_),
    .A(_2433_),
    .B(_2445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3098_ (.A(_2437_),
    .B(_2446_),
    .Y(_2447_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3099_ (.B1(net816),
    .VDD(VPWR),
    .Y(_2448_),
    .VSS(VGND),
    .A1(net901),
    .A2(net1002));
 sg13g2_a21oi_1 _3100_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(net1002),
    .Y(_0005_),
    .B1(_2448_));
 sg13g2_nor2b_2 _3101_ (.A(net1132),
    .B_N(\falu_i.falutop.i2c_inst.counter[1] ),
    .Y(_0343_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3102_ (.Y(_0344_),
    .A(_2433_),
    .B(net1046),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3103_ (.A(net1014),
    .B(_0344_),
    .Y(_0345_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3104_ (.B1(net820),
    .VDD(VPWR),
    .Y(_0346_),
    .VSS(VGND),
    .A1(net972),
    .A2(_0345_));
 sg13g2_a21oi_1 _3105_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net801),
    .A2(_0345_),
    .Y(_0006_),
    .B1(_0346_));
 sg13g2_nor2_1 _3106_ (.A(_2434_),
    .B(net1014),
    .Y(_0347_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3107_ (.B1(net823),
    .VDD(VPWR),
    .Y(_0348_),
    .VSS(VGND),
    .A1(net992),
    .A2(_0347_));
 sg13g2_a21oi_1 _3108_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net801),
    .A2(_0347_),
    .Y(_0007_),
    .B1(_0348_));
 sg13g2_nor2_1 _3109_ (.A(net985),
    .B(_2154_),
    .Y(_0349_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3110_ (.Y(_0350_),
    .B(_0349_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\falu_i.falutop.i2c_inst.counter[4] ));
 sg13g2_nor2_1 _3111_ (.A(_2439_),
    .B(net987),
    .Y(_0351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3112_ (.B1(net817),
    .VDD(VPWR),
    .Y(_0352_),
    .VSS(VGND),
    .A1(net881),
    .A2(net988));
 sg13g2_a21oi_1 _3113_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(net988),
    .Y(_0008_),
    .B1(_0352_));
 sg13g2_nor2_1 _3114_ (.A(_2446_),
    .B(net987),
    .Y(_0353_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3115_ (.B1(net804),
    .VDD(VPWR),
    .Y(_0354_),
    .VSS(VGND),
    .A1(net869),
    .A2(_0353_));
 sg13g2_a21oi_1 _3116_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0353_),
    .Y(_0009_),
    .B1(_0354_));
 sg13g2_nor2_1 _3117_ (.A(_0344_),
    .B(net987),
    .Y(_0355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3118_ (.B1(net804),
    .VDD(VPWR),
    .Y(_0356_),
    .VSS(VGND),
    .A1(net850),
    .A2(_0355_));
 sg13g2_a21oi_1 _3119_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0355_),
    .Y(_0010_),
    .B1(_0356_));
 sg13g2_nor2_1 _3120_ (.A(_2434_),
    .B(net987),
    .Y(_0357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3121_ (.B1(net804),
    .VDD(VPWR),
    .Y(_0358_),
    .VSS(VGND),
    .A1(net871),
    .A2(_0357_));
 sg13g2_a21oi_1 _3122_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0357_),
    .Y(_0011_),
    .B1(_0358_));
 sg13g2_nor2b_2 _3123_ (.A(net1016),
    .B_N(\falu_i.falutop.i2c_inst.counter[3] ),
    .Y(_0359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3124_ (.Y(_0360_),
    .A(_2154_),
    .B(net1017),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3125_ (.A(_2439_),
    .B(_0360_),
    .Y(_0361_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3126_ (.B1(net804),
    .VDD(VPWR),
    .Y(_0362_),
    .VSS(VGND),
    .A1(net873),
    .A2(_0361_));
 sg13g2_a21oi_1 _3127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0361_),
    .Y(_0012_),
    .B1(_0362_));
 sg13g2_nor2_1 _3128_ (.A(_2446_),
    .B(_0360_),
    .Y(_0363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3129_ (.B1(net820),
    .VDD(VPWR),
    .Y(_0364_),
    .VSS(VGND),
    .A1(net899),
    .A2(_0363_));
 sg13g2_a21oi_1 _3130_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0363_),
    .Y(_0013_),
    .B1(_0364_));
 sg13g2_nor2_1 _3131_ (.A(_0344_),
    .B(_0360_),
    .Y(_0365_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3132_ (.B1(net816),
    .VDD(VPWR),
    .Y(_0366_),
    .VSS(VGND),
    .A1(net945),
    .A2(_0365_));
 sg13g2_a21oi_1 _3133_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0365_),
    .Y(_0014_),
    .B1(_0366_));
 sg13g2_nor2_1 _3134_ (.A(_2434_),
    .B(_0360_),
    .Y(_0367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3135_ (.B1(net816),
    .VDD(VPWR),
    .Y(_0368_),
    .VSS(VGND),
    .A1(net858),
    .A2(_0367_));
 sg13g2_a21oi_1 _3136_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0367_),
    .Y(_0015_),
    .B1(_0368_));
 sg13g2_nand2_2 _3137_ (.Y(_0369_),
    .A(net1006),
    .B(_0359_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3138_ (.A(_2439_),
    .B(net1007),
    .Y(_0370_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3139_ (.B1(net816),
    .VDD(VPWR),
    .Y(_0371_),
    .VSS(VGND),
    .A1(net926),
    .A2(_0370_));
 sg13g2_a21oi_1 _3140_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0370_),
    .Y(_0016_),
    .B1(_0371_));
 sg13g2_nor2_1 _3141_ (.A(_2446_),
    .B(net1007),
    .Y(_0372_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3142_ (.B1(net816),
    .VDD(VPWR),
    .Y(_0373_),
    .VSS(VGND),
    .A1(net894),
    .A2(_0372_));
 sg13g2_a21oi_1 _3143_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0372_),
    .Y(_0017_),
    .B1(_0373_));
 sg13g2_nor2_1 _3144_ (.A(_0344_),
    .B(net1007),
    .Y(_0374_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3145_ (.B1(net804),
    .VDD(VPWR),
    .Y(_0375_),
    .VSS(VGND),
    .A1(net861),
    .A2(_0374_));
 sg13g2_a21oi_1 _3146_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0374_),
    .Y(_0018_),
    .B1(_0375_));
 sg13g2_nor2_1 _3147_ (.A(_2434_),
    .B(net1007),
    .Y(_0376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3148_ (.B1(net804),
    .VDD(VPWR),
    .Y(_0377_),
    .VSS(VGND),
    .A1(net908),
    .A2(_0376_));
 sg13g2_a21oi_1 _3149_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net802),
    .A2(_0376_),
    .Y(_0019_),
    .B1(_0377_));
 sg13g2_nor2_1 _3150_ (.A(_2431_),
    .B(_2439_),
    .Y(_0378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3151_ (.B1(net820),
    .VDD(VPWR),
    .Y(_0379_),
    .VSS(VGND),
    .A1(net1070),
    .A2(_0378_));
 sg13g2_a21oi_1 _3152_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net800),
    .A2(_0378_),
    .Y(_0020_),
    .B1(_0379_));
 sg13g2_nor2_1 _3153_ (.A(_2431_),
    .B(_2446_),
    .Y(_0380_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3154_ (.B1(net821),
    .VDD(VPWR),
    .Y(_0381_),
    .VSS(VGND),
    .A1(net912),
    .A2(_0380_));
 sg13g2_a21oi_1 _3155_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net801),
    .A2(_0380_),
    .Y(_0021_),
    .B1(_0381_));
 sg13g2_nor2_1 _3156_ (.A(_2431_),
    .B(_0344_),
    .Y(_0382_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3157_ (.B1(net820),
    .VDD(VPWR),
    .Y(_0383_),
    .VSS(VGND),
    .A1(net1044),
    .A2(_0382_));
 sg13g2_a21oi_1 _3158_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net801),
    .A2(_0382_),
    .Y(_0022_),
    .B1(_0383_));
 sg13g2_and2_1 _3159_ (.A(net807),
    .B(net373),
    .X(_0023_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3160_ (.A(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .B(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .C(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .Y(_0384_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3161_ (.A(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .B(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .C(\ppwm_i.u_ppwm.u_pwm.counter[5] ),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .Y(_0385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3162_ (.B(_2274_),
    .C(_0384_),
    .A(_2273_),
    .Y(_0386_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0385_));
 sg13g2_o21ai_1 _3163_ (.B1(net811),
    .VDD(VPWR),
    .Y(_0387_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[0] ),
    .A2(net681));
 sg13g2_a21oi_1 _3164_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2288_),
    .A2(net681),
    .Y(_0024_),
    .B1(_0387_));
 sg13g2_o21ai_1 _3165_ (.B1(net807),
    .VDD(VPWR),
    .Y(_0388_),
    .VSS(VGND),
    .A1(net785),
    .A2(net681));
 sg13g2_a21oi_1 _3166_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2287_),
    .A2(net681),
    .Y(_0025_),
    .B1(_0388_));
 sg13g2_o21ai_1 _3167_ (.B1(net808),
    .VDD(VPWR),
    .Y(_0389_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[2] ),
    .A2(net681));
 sg13g2_a21oi_1 _3168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2286_),
    .A2(net681),
    .Y(_0026_),
    .B1(_0389_));
 sg13g2_o21ai_1 _3169_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0390_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[3] ),
    .A2(net681));
 sg13g2_a21oi_1 _3170_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2285_),
    .A2(net683),
    .Y(_0027_),
    .B1(_0390_));
 sg13g2_o21ai_1 _3171_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0391_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A2(net683));
 sg13g2_a21oi_1 _3172_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2284_),
    .A2(net681),
    .Y(_0028_),
    .B1(_0391_));
 sg13g2_o21ai_1 _3173_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0392_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[5] ),
    .A2(net682));
 sg13g2_a21oi_1 _3174_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2283_),
    .A2(net682),
    .Y(_0029_),
    .B1(_0392_));
 sg13g2_o21ai_1 _3175_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0393_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[6] ),
    .A2(net682));
 sg13g2_a21oi_1 _3176_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2282_),
    .A2(net682),
    .Y(_0030_),
    .B1(_0393_));
 sg13g2_o21ai_1 _3177_ (.B1(net813),
    .VDD(VPWR),
    .Y(_0394_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[7] ),
    .A2(net682));
 sg13g2_a21oi_1 _3178_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2281_),
    .A2(net683),
    .Y(_0031_),
    .B1(_0394_));
 sg13g2_o21ai_1 _3179_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0395_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .A2(net682));
 sg13g2_a21oi_1 _3180_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2280_),
    .A2(net682),
    .Y(_0032_),
    .B1(_0395_));
 sg13g2_o21ai_1 _3181_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0396_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[9] ),
    .A2(net682));
 sg13g2_a21oi_1 _3182_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2279_),
    .A2(net683),
    .Y(_0033_),
    .B1(_0396_));
 sg13g2_nand2_1 _3183_ (.Y(_0397_),
    .A(net512),
    .B(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3184_ (.B(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .C(net1010),
    .A(net512),
    .Y(_0398_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2155_));
 sg13g2_nor4_1 _3185_ (.A(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .B(\ppwm_i.u_ppwm.u_mem.bit_count[1] ),
    .C(net378),
    .D(_0398_),
    .Y(_0399_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3186_ (.A(net1111),
    .B(_0399_),
    .X(_0400_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3187_ (.B1(net807),
    .VDD(VPWR),
    .Y(_0401_),
    .VSS(VGND),
    .A1(net1111),
    .A2(_0399_));
 sg13g2_nor2_1 _3188_ (.A(_0400_),
    .B(net1112),
    .Y(_0034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3189_ (.A(net1117),
    .B(_0400_),
    .X(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3190_ (.B1(net808),
    .VDD(VPWR),
    .Y(_0403_),
    .VSS(VGND),
    .A1(net1117),
    .A2(_0400_));
 sg13g2_nor2_1 _3191_ (.A(_0402_),
    .B(net1118),
    .Y(_0035_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3192_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0404_),
    .B(_0402_),
    .A(net1049));
 sg13g2_nand2_1 _3193_ (.Y(_0405_),
    .A(net1049),
    .B(_0402_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3194_ (.X(_0036_),
    .A(net809),
    .B(_0404_),
    .C(net1050),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3195_ (.Y(_0406_),
    .A(net863),
    .B(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3196_ (.B(net1049),
    .C(_0402_),
    .A(net863),
    .Y(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3197_ (.Y(_0408_),
    .A(net809),
    .B(_0407_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3198_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2278_),
    .A2(net1050),
    .Y(_0037_),
    .B1(_0408_));
 sg13g2_or2_1 _3199_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0409_),
    .B(_0407_),
    .A(_2277_));
 sg13g2_nand2_1 _3200_ (.Y(_0410_),
    .A(net809),
    .B(_0409_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3201_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2277_),
    .A2(_0407_),
    .Y(_0038_),
    .B1(_0410_));
 sg13g2_nand2_2 _3202_ (.Y(_0411_),
    .A(net1060),
    .B(net1090),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3203_ (.A(_0407_),
    .B(_0411_),
    .Y(_0412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3204_ (.B1(net809),
    .VDD(VPWR),
    .Y(_0413_),
    .VSS(VGND),
    .A1(_0407_),
    .A2(_0411_));
 sg13g2_a21oi_1 _3205_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2276_),
    .A2(_0409_),
    .Y(_0039_),
    .B1(_0413_));
 sg13g2_nor2_1 _3206_ (.A(net1066),
    .B(_0412_),
    .Y(_0414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3207_ (.A(_2275_),
    .B(_0407_),
    .C(_0411_),
    .Y(_0415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3208_ (.A(net796),
    .B(net1067),
    .C(_0415_),
    .Y(_0040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3209_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0416_),
    .B(_0415_),
    .A(net1177));
 sg13g2_nand2_1 _3210_ (.Y(_0417_),
    .A(net1177),
    .B(_0415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3211_ (.X(_0041_),
    .A(net809),
    .B(_0416_),
    .C(_0417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3212_ (.B(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .C(_0415_),
    .A(net1094),
    .Y(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3213_ (.Y(_0419_),
    .A(net809),
    .B(_0418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3214_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2274_),
    .A2(_0417_),
    .Y(_0042_),
    .B1(_0419_));
 sg13g2_o21ai_1 _3215_ (.B1(net809),
    .VDD(VPWR),
    .Y(_0420_),
    .VSS(VGND),
    .A1(_2273_),
    .A2(_0418_));
 sg13g2_a21oi_1 _3216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2273_),
    .A2(_0418_),
    .Y(_0043_),
    .B1(_0420_));
 sg13g2_nand3_1 _3217_ (.B(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .C(net809),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .Y(_0421_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3218_ (.B(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .C(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .A(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .Y(_0422_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(\ppwm_i.u_ppwm.u_pwm.counter[6] ));
 sg13g2_nor4_1 _3219_ (.A(net864),
    .B(_0411_),
    .C(_0421_),
    .D(_0422_),
    .Y(_0044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3220_ (.Y(_0423_),
    .A(net1039),
    .B(net1096),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3221_ (.A(net795),
    .B(_0423_),
    .Y(_0045_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3222_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.period_start ),
    .A2(\ppwm_i.u_ppwm.global_counter[0] ),
    .Y(_0424_),
    .B1(net942));
 sg13g2_nand3_1 _3223_ (.B(net942),
    .C(\ppwm_i.u_ppwm.global_counter[0] ),
    .A(\ppwm_i.u_ppwm.period_start ),
    .Y(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3224_ (.Y(_0426_),
    .A(net812),
    .B(_0425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3225_ (.A(net943),
    .B(_0426_),
    .Y(_0046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3226_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0427_),
    .B(_0425_),
    .A(_2272_));
 sg13g2_nand2_1 _3227_ (.Y(_0428_),
    .A(net812),
    .B(_0427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3228_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2272_),
    .A2(_0425_),
    .Y(_0047_),
    .B1(_0428_));
 sg13g2_and2_1 _3229_ (.A(_2271_),
    .B(_0427_),
    .X(_0429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3230_ (.A(_2271_),
    .B(_0427_),
    .Y(_0430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3231_ (.A(net795),
    .B(_0429_),
    .C(_0430_),
    .Y(_0048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _3232_ (.A(_2270_),
    .B(_2271_),
    .C(_0427_),
    .Y(_0431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3233_ (.B1(net812),
    .VDD(VPWR),
    .Y(_0432_),
    .VSS(VGND),
    .A1(net1107),
    .A2(_0430_));
 sg13g2_nor2_1 _3234_ (.A(_0431_),
    .B(net1108),
    .Y(_0049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3235_ (.Y(_0433_),
    .A(net1145),
    .B(_0431_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3236_ (.B1(net813),
    .VDD(VPWR),
    .Y(_0434_),
    .VSS(VGND),
    .A1(net1145),
    .A2(_0431_));
 sg13g2_nor2b_1 _3237_ (.A(net1146),
    .B_N(_0433_),
    .Y(_0050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3238_ (.A(_2269_),
    .B(_0433_),
    .Y(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3239_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2269_),
    .A2(_0433_),
    .Y(_0436_),
    .B1(net795));
 sg13g2_nor2b_1 _3240_ (.A(_0435_),
    .B_N(net1185),
    .Y(_0051_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3241_ (.Y(_0437_),
    .A(net1092),
    .B(_0435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3242_ (.A(net796),
    .B(net1093),
    .Y(_0052_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3243_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[7] ),
    .A2(_0435_),
    .Y(_0438_),
    .B1(net553));
 sg13g2_nor4_1 _3244_ (.A(_2267_),
    .B(_2268_),
    .C(_2269_),
    .D(_0433_),
    .Y(_0439_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3245_ (.A(net795),
    .B(net554),
    .C(_0439_),
    .Y(_0053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3246_ (.A(net1139),
    .B(_0439_),
    .X(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3247_ (.B1(net812),
    .VDD(VPWR),
    .Y(_0441_),
    .VSS(VGND),
    .A1(net1139),
    .A2(_0439_));
 sg13g2_nor2_1 _3248_ (.A(_0440_),
    .B(net1140),
    .Y(_0054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3249_ (.Y(_0442_),
    .A(net1120),
    .B(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3250_ (.A(net795),
    .B(net1121),
    .Y(_0055_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3251_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[10] ),
    .A2(_0440_),
    .Y(_0443_),
    .B1(net954));
 sg13g2_and3_1 _3252_ (.X(_0444_),
    .A(net954),
    .B(net1120),
    .C(_0440_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3253_ (.A(net795),
    .B(net955),
    .C(_0444_),
    .Y(_0056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3254_ (.A(net1134),
    .B(_0444_),
    .X(_0445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3255_ (.B1(net812),
    .VDD(VPWR),
    .Y(_0446_),
    .VSS(VGND),
    .A1(net1134),
    .A2(_0444_));
 sg13g2_nor2_1 _3256_ (.A(_0445_),
    .B(_0446_),
    .Y(_0057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3257_ (.Y(_0447_),
    .A(net1129),
    .B(_0445_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3258_ (.A(net796),
    .B(net1130),
    .Y(_0058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3259_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[13] ),
    .A2(_0445_),
    .Y(_0448_),
    .B1(net974));
 sg13g2_nand3_1 _3260_ (.B(net1129),
    .C(_0445_),
    .A(net974),
    .Y(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3261_ (.Y(_0450_),
    .A(net812),
    .B(_0449_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3262_ (.A(net975),
    .B(_0450_),
    .Y(_0059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3263_ (.A(_2262_),
    .B(_0449_),
    .X(_0451_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3264_ (.A(_2262_),
    .B(_0449_),
    .Y(_0452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3265_ (.A(net796),
    .B(_0451_),
    .C(_0452_),
    .Y(_0060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3266_ (.Y(_0453_),
    .A(net1125),
    .B(_0452_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3267_ (.A(net796),
    .B(net1126),
    .Y(_0061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3268_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[16] ),
    .A2(_0452_),
    .Y(_0454_),
    .B1(net989));
 sg13g2_nand3_1 _3269_ (.B(\ppwm_i.u_ppwm.global_counter[16] ),
    .C(_0452_),
    .A(net989),
    .Y(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3270_ (.Y(_0456_),
    .A(net812),
    .B(_0455_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3271_ (.A(net990),
    .B(_0456_),
    .Y(_0062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3272_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0457_),
    .B(_0455_),
    .A(_2259_));
 sg13g2_nand2_1 _3273_ (.Y(_0458_),
    .A(net813),
    .B(_0457_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3274_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2259_),
    .A2(_0455_),
    .Y(_0063_),
    .B1(_0458_));
 sg13g2_o21ai_1 _3275_ (.B1(net812),
    .VDD(VPWR),
    .Y(_0459_),
    .VSS(VGND),
    .A1(_2258_),
    .A2(_0457_));
 sg13g2_a21oi_1 _3276_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2258_),
    .A2(_0457_),
    .Y(_0064_),
    .B1(_0459_));
 sg13g2_nand2b_1 _3277_ (.Y(_0460_),
    .B(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ),
    .A_N(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3278_ (.B1(_0460_),
    .VDD(VPWR),
    .Y(_0461_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .A2(_2288_));
 sg13g2_a22oi_1 _3279_ (.Y(_0462_),
    .B1(_2287_),
    .B2(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .A2(_2286_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3280_ (.A(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .B(_2286_),
    .Y(_0463_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3281_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0462_),
    .C1(_0463_),
    .B1(_0461_),
    .A1(_2278_),
    .Y(_0464_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[3] ));
 sg13g2_a221oi_1 _3282_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .C1(_0464_),
    .B1(_2285_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .Y(_0465_),
    .A2(_2284_));
 sg13g2_a21oi_1 _3283_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2277_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[4] ),
    .Y(_0466_),
    .B1(_0465_));
 sg13g2_a21o_1 _3284_ (.A2(_2283_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[5] ),
    .B1(_0466_),
    .X(_0467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3285_ (.Y(_0468_),
    .B1(\ppwm_i.u_ppwm.u_pwm.cmp_value[5] ),
    .B2(_2276_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ),
    .A1(_2275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3286_ (.Y(_0469_),
    .B1(_0467_),
    .B2(_0468_),
    .A2(_2281_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3287_ (.B1(_0469_),
    .VDD(VPWR),
    .Y(_0470_),
    .VSS(VGND),
    .A1(_2275_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ));
 sg13g2_o21ai_1 _3288_ (.B1(_0470_),
    .VDD(VPWR),
    .Y(_0471_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .A2(_2281_));
 sg13g2_a21oi_1 _3289_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2274_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[8] ),
    .Y(_0472_),
    .B1(_0471_));
 sg13g2_a221oi_1 _3290_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .C1(_0472_),
    .B1(_2280_),
    .A1(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .Y(_0473_),
    .A2(_2279_));
 sg13g2_a21oi_1 _3291_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2273_),
    .A2(\ppwm_i.u_ppwm.u_pwm.cmp_value[9] ),
    .Y(_0474_),
    .B1(_0473_));
 sg13g2_o21ai_1 _3292_ (.B1(net810),
    .VDD(VPWR),
    .Y(_0475_),
    .VSS(VGND),
    .A1(net376),
    .A2(_0474_));
 sg13g2_a21oi_1 _3293_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net376),
    .A2(_0474_),
    .Y(_0065_),
    .B1(_0475_));
 sg13g2_nand2_1 _3294_ (.Y(_0476_),
    .A(net793),
    .B(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3295_ (.Y(_0477_),
    .A(_2257_),
    .B(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3296_ (.Y(_0478_),
    .B(_2360_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2344_));
 sg13g2_or2_1 _3297_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0479_),
    .B(_0478_),
    .A(_2329_));
 sg13g2_a21oi_1 _3298_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2253_),
    .A2(net793),
    .Y(_0480_),
    .B1(_0479_));
 sg13g2_o21ai_1 _3299_ (.B1(_0480_),
    .VDD(VPWR),
    .Y(_0481_),
    .VSS(VGND),
    .A1(_2253_),
    .A2(_0477_));
 sg13g2_nor2_2 _3300_ (.A(_2330_),
    .B(_0478_),
    .Y(_0482_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3301_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0477_),
    .C1(_2255_),
    .B1(_0482_),
    .A1(_2257_),
    .Y(_0483_),
    .A2(_0478_));
 sg13g2_a221oi_1 _3302_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0483_),
    .C1(net799),
    .B1(net1163),
    .A1(_2255_),
    .Y(_0066_),
    .A2(_2257_));
 sg13g2_a21oi_1 _3303_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2307_),
    .A2(_2310_),
    .Y(_0484_),
    .B1(net1162));
 sg13g2_xnor2_1 _3304_ (.Y(_0485_),
    .A(net791),
    .B(_2418_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3305_ (.A(_0476_),
    .B(_0485_),
    .Y(_0486_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3306_ (.Y(_0487_),
    .A(_0476_),
    .B(_0485_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3307_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1162),
    .A2(_0487_),
    .Y(_0488_),
    .B1(_0484_));
 sg13g2_o21ai_1 _3308_ (.B1(_0478_),
    .VDD(VPWR),
    .Y(_0489_),
    .VSS(VGND),
    .A1(net700),
    .A2(net696));
 sg13g2_nand2b_1 _3309_ (.Y(_0490_),
    .B(_0489_),
    .A_N(_2422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3310_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0482_),
    .A2(_0487_),
    .Y(_0491_),
    .B1(_0490_));
 sg13g2_o21ai_1 _3311_ (.B1(_0491_),
    .VDD(VPWR),
    .Y(_0492_),
    .VSS(VGND),
    .A1(_0479_),
    .A2(_0488_));
 sg13g2_nor2_1 _3312_ (.A(net419),
    .B(net799),
    .Y(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3313_ (.Y(_0494_),
    .A(net791),
    .B(_0493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3314_ (.Y(_0067_),
    .A(_0492_),
    .B(_0494_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3315_ (.Y(_0495_),
    .A(net788),
    .B(net701),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3316_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net791),
    .A2(_2418_),
    .Y(_0496_),
    .B1(_0486_));
 sg13g2_nand2_1 _3317_ (.Y(_0497_),
    .A(net788),
    .B(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3318_ (.Y(_0498_),
    .A(net788),
    .B(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3319_ (.Y(_0499_),
    .A(_0496_),
    .B(_0498_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3320_ (.A(net1162),
    .B(_0495_),
    .Y(_0500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3321_ (.A(_0479_),
    .B(_0500_),
    .Y(_0501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3322_ (.B1(_0501_),
    .VDD(VPWR),
    .Y(_0502_),
    .VSS(VGND),
    .A1(_2253_),
    .A2(_0499_));
 sg13g2_a221oi_1 _3323_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0482_),
    .C1(_2422_),
    .B1(_0499_),
    .A1(_0478_),
    .Y(_0503_),
    .A2(_0495_));
 sg13g2_a22oi_1 _3324_ (.Y(_0504_),
    .B1(_0502_),
    .B2(_0503_),
    .A2(_0493_),
    .A1(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3325_ (.VDD(VPWR),
    .Y(_0068_),
    .A(_0504_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3326_ (.B1(_2254_),
    .VDD(VPWR),
    .Y(_0505_),
    .VSS(VGND),
    .A1(net708),
    .A2(_2307_));
 sg13g2_nand2_1 _3327_ (.Y(_0506_),
    .A(_2308_),
    .B(_0505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3328_ (.A(_2254_),
    .B(_2367_),
    .Y(_0507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3329_ (.A(_2373_),
    .B(_0507_),
    .Y(_0508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3330_ (.B1(_0497_),
    .VDD(VPWR),
    .Y(_0509_),
    .VSS(VGND),
    .A1(_0496_),
    .A2(_0498_));
 sg13g2_xor2_1 _3331_ (.B(_0509_),
    .A(_0508_),
    .X(_0510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3332_ (.A(net1162),
    .B(_0506_),
    .Y(_0511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3333_ (.A(_0479_),
    .B(_0511_),
    .Y(_0512_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3334_ (.B1(_0512_),
    .VDD(VPWR),
    .Y(_0513_),
    .VSS(VGND),
    .A1(_2253_),
    .A2(_0510_));
 sg13g2_a221oi_1 _3335_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0482_),
    .C1(_2422_),
    .B1(_0510_),
    .A1(_0478_),
    .Y(_0514_),
    .A2(_0506_));
 sg13g2_a22oi_1 _3336_ (.Y(_0515_),
    .B1(_0513_),
    .B2(_0514_),
    .A2(_0493_),
    .A1(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3337_ (.VDD(VPWR),
    .Y(_0069_),
    .A(_0515_),
    .VSS(VGND));
 sg13g2_nand4_1 _3338_ (.B(_2330_),
    .C(_2344_),
    .A(net419),
    .Y(_0516_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2360_));
 sg13g2_nand2_1 _3339_ (.Y(_0517_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .B(_2243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3340_ (.A(net782),
    .B(_2244_),
    .Y(_0518_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3341_ (.Y(_0519_),
    .A(_2242_),
    .B(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3342_ (.A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .B_N(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .Y(_0520_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3343_ (.A(_2242_),
    .B(net784),
    .Y(_0521_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3344_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0520_),
    .C1(_0521_),
    .B1(_0519_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .Y(_0522_),
    .A2(_2250_));
 sg13g2_a221oi_1 _3345_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2241_),
    .C1(_0522_),
    .B1(\ppwm_i.u_ppwm.pwm_value[2] ),
    .A1(_2240_),
    .Y(_0523_),
    .A2(\ppwm_i.u_ppwm.pwm_value[3] ));
 sg13g2_a221oi_1 _3346_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .C1(_0523_),
    .B1(_2249_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .Y(_0524_),
    .A2(_2248_));
 sg13g2_a221oi_1 _3347_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2239_),
    .C1(_0524_),
    .B1(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A1(_2238_),
    .Y(_0525_),
    .A2(\ppwm_i.u_ppwm.pwm_value[5] ));
 sg13g2_a221oi_1 _3348_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .C1(_0525_),
    .B1(_2247_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .Y(_0526_),
    .A2(_2246_));
 sg13g2_a221oi_1 _3349_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2237_),
    .C1(_0526_),
    .B1(\ppwm_i.u_ppwm.pwm_value[6] ),
    .A1(_2236_),
    .Y(_0527_),
    .A2(\ppwm_i.u_ppwm.pwm_value[7] ));
 sg13g2_a221oi_1 _3350_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .C1(_0527_),
    .B1(_2245_),
    .A1(net782),
    .Y(_0528_),
    .A2(_2244_));
 sg13g2_o21ai_1 _3351_ (.B1(_0517_),
    .VDD(VPWR),
    .Y(_0529_),
    .VSS(VGND),
    .A1(_0518_),
    .A2(_0528_));
 sg13g2_nor2_1 _3352_ (.A(net612),
    .B(_2419_),
    .Y(_0530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3353_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2235_),
    .A2(\ppwm_i.u_ppwm.pwm_value[9] ),
    .Y(_0531_),
    .B1(net591));
 sg13g2_nand3_1 _3354_ (.B(net581),
    .C(_0531_),
    .A(_0529_),
    .Y(_0532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3355_ (.A(\ppwm_i.u_ppwm.pwm_value[7] ),
    .B(_2268_),
    .Y(_0533_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3356_ (.Y(_0534_),
    .B(\ppwm_i.u_ppwm.global_counter[1] ),
    .A_N(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3357_ (.B(_0534_),
    .C(\ppwm_i.u_ppwm.pwm_value[0] ),
    .Y(_0535_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\ppwm_i.u_ppwm.global_counter[0] ));
 sg13g2_nand2b_1 _3358_ (.Y(_0536_),
    .B(net784),
    .A_N(\ppwm_i.u_ppwm.global_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3359_ (.Y(_0537_),
    .B1(_0535_),
    .B2(_0536_),
    .A2(\ppwm_i.u_ppwm.global_counter[2] ),
    .A1(_2250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3360_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.pwm_value[2] ),
    .C1(_0537_),
    .B1(_2272_),
    .A1(\ppwm_i.u_ppwm.pwm_value[3] ),
    .Y(_0538_),
    .A2(_2271_));
 sg13g2_a221oi_1 _3361_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2249_),
    .C1(_0538_),
    .B1(\ppwm_i.u_ppwm.global_counter[3] ),
    .A1(_2248_),
    .Y(_0539_),
    .A2(\ppwm_i.u_ppwm.global_counter[4] ));
 sg13g2_a21oi_1 _3362_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A2(_2270_),
    .Y(_0540_),
    .B1(_0539_));
 sg13g2_o21ai_1 _3363_ (.B1(_0540_),
    .VDD(VPWR),
    .Y(_0541_),
    .VSS(VGND),
    .A1(_2247_),
    .A2(\ppwm_i.u_ppwm.global_counter[5] ));
 sg13g2_a22oi_1 _3364_ (.Y(_0542_),
    .B1(\ppwm_i.u_ppwm.global_counter[5] ),
    .B2(_2247_),
    .A2(\ppwm_i.u_ppwm.global_counter[6] ),
    .A1(_2246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3365_ (.Y(_0543_),
    .B1(_0541_),
    .B2(_0542_),
    .A2(_2269_),
    .A1(\ppwm_i.u_ppwm.pwm_value[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3366_ (.Y(_0544_),
    .B1(_2268_),
    .B2(\ppwm_i.u_ppwm.pwm_value[7] ),
    .A2(_2267_),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3367_ (.B1(_0544_),
    .VDD(VPWR),
    .Y(_0545_),
    .VSS(VGND),
    .A1(_0533_),
    .A2(_0543_));
 sg13g2_o21ai_1 _3368_ (.B1(_0545_),
    .VDD(VPWR),
    .Y(_0546_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .A2(_2267_));
 sg13g2_o21ai_1 _3369_ (.B1(_0546_),
    .VDD(VPWR),
    .Y(_0547_),
    .VSS(VGND),
    .A1(_2243_),
    .A2(\ppwm_i.u_ppwm.global_counter[9] ));
 sg13g2_nor2_1 _3370_ (.A(_2243_),
    .B(net596),
    .Y(_0548_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3371_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2243_),
    .A2(\ppwm_i.u_ppwm.global_counter[9] ),
    .Y(_0549_),
    .B1(net591));
 sg13g2_nand2_1 _3372_ (.Y(_0550_),
    .A(_2237_),
    .B(\ppwm_i.u_ppwm.global_counter[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3373_ (.A(_2238_),
    .B(\ppwm_i.u_ppwm.global_counter[5] ),
    .Y(_0551_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3374_ (.Y(_0552_),
    .A(_2240_),
    .B(\ppwm_i.u_ppwm.global_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3375_ (.Y(_0553_),
    .B(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .A_N(\ppwm_i.u_ppwm.global_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3376_ (.B1(_0553_),
    .VDD(VPWR),
    .Y(_0554_),
    .VSS(VGND),
    .A1(_2242_),
    .A2(\ppwm_i.u_ppwm.global_counter[1] ));
 sg13g2_a22oi_1 _3377_ (.Y(_0555_),
    .B1(\ppwm_i.u_ppwm.global_counter[1] ),
    .B2(_2242_),
    .A2(\ppwm_i.u_ppwm.global_counter[2] ),
    .A1(_2241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3378_ (.Y(_0556_),
    .B1(_0554_),
    .B2(_0555_),
    .A2(_2271_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3379_ (.B1(_0556_),
    .VDD(VPWR),
    .Y(_0557_),
    .VSS(VGND),
    .A1(_2241_),
    .A2(\ppwm_i.u_ppwm.global_counter[2] ));
 sg13g2_a22oi_1 _3380_ (.Y(_0558_),
    .B1(_0552_),
    .B2(_0557_),
    .A2(_2270_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3381_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2239_),
    .C1(_0558_),
    .B1(\ppwm_i.u_ppwm.global_counter[4] ),
    .A1(_2238_),
    .Y(_0559_),
    .A2(\ppwm_i.u_ppwm.global_counter[5] ));
 sg13g2_o21ai_1 _3382_ (.B1(_0550_),
    .VDD(VPWR),
    .Y(_0560_),
    .VSS(VGND),
    .A1(_0551_),
    .A2(_0559_));
 sg13g2_a22oi_1 _3383_ (.Y(_0561_),
    .B1(_2269_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .A2(_2268_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3384_ (.Y(_0562_),
    .B1(_0560_),
    .B2(_0561_),
    .A2(\ppwm_i.u_ppwm.global_counter[7] ),
    .A1(_2236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3385_ (.A(_2235_),
    .B(\ppwm_i.u_ppwm.global_counter[9] ),
    .Y(_0563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3386_ (.B(\ppwm_i.u_ppwm.global_counter[8] ),
    .A(net782),
    .X(_0564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3387_ (.A(_0562_),
    .B(_0563_),
    .C(_0564_),
    .Y(_0565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3388_ (.Y(_0566_),
    .A(_2235_),
    .B(\ppwm_i.u_ppwm.global_counter[9] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3389_ (.A(net782),
    .B(_2267_),
    .C(_0563_),
    .Y(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3390_ (.Y(_0568_),
    .B(net592),
    .A_N(_0567_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3391_ (.A(_0565_),
    .B(_0568_),
    .Y(_0569_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3392_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0569_),
    .C1(net610),
    .B1(_0566_),
    .A1(_0547_),
    .Y(_0570_),
    .A2(_0549_));
 sg13g2_nor2b_1 _3393_ (.A(\ppwm_i.u_ppwm.global_counter[10] ),
    .B_N(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .Y(_0571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3394_ (.B1(_0571_),
    .VDD(VPWR),
    .Y(_0572_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .A2(_2266_));
 sg13g2_a22oi_1 _3395_ (.Y(_0573_),
    .B1(_2266_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .A2(_2265_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3396_ (.Y(_0574_),
    .B1(_0572_),
    .B2(_0573_),
    .A2(\ppwm_i.u_ppwm.global_counter[12] ),
    .A1(_2241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3397_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .A2(_2264_),
    .Y(_0575_),
    .B1(_0574_));
 sg13g2_a221oi_1 _3398_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2240_),
    .C1(_0575_),
    .B1(\ppwm_i.u_ppwm.global_counter[13] ),
    .A1(_2239_),
    .Y(_0576_),
    .A2(\ppwm_i.u_ppwm.global_counter[14] ));
 sg13g2_a221oi_1 _3399_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .C1(_0576_),
    .B1(_2263_),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .Y(_0577_),
    .A2(_2262_));
 sg13g2_a221oi_1 _3400_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2238_),
    .C1(_0577_),
    .B1(\ppwm_i.u_ppwm.global_counter[15] ),
    .A1(_2237_),
    .Y(_0578_),
    .A2(\ppwm_i.u_ppwm.global_counter[16] ));
 sg13g2_a21oi_1 _3401_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .A2(_2261_),
    .Y(_0579_),
    .B1(_0578_));
 sg13g2_a21o_1 _3402_ (.A2(\ppwm_i.u_ppwm.global_counter[17] ),
    .A1(_2236_),
    .B1(_0579_),
    .X(_0580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3403_ (.Y(_0581_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .B(_2258_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3404_ (.Y(_0582_),
    .B(\ppwm_i.u_ppwm.global_counter[18] ),
    .A_N(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3405_ (.Y(_0583_),
    .B1(_2260_),
    .B2(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .A2(_2259_),
    .A1(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3406_ (.B(_0581_),
    .C(_0582_),
    .A(_0580_),
    .Y(_0584_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0583_));
 sg13g2_nand3b_1 _3407_ (.B(\ppwm_i.u_ppwm.global_counter[18] ),
    .C(_0581_),
    .Y(_0585_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net782));
 sg13g2_nand2_1 _3408_ (.Y(_0586_),
    .A(_2258_),
    .B(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3409_ (.Y(_0587_),
    .A(_2235_),
    .B(\ppwm_i.u_ppwm.global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3410_ (.B(_0584_),
    .C(_0585_),
    .A(net591),
    .Y(_0588_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0587_));
 sg13g2_a21oi_1 _3411_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2243_),
    .A2(\ppwm_i.u_ppwm.global_counter[19] ),
    .Y(_0589_),
    .B1(net591));
 sg13g2_nor2_1 _3412_ (.A(net784),
    .B(_2266_),
    .Y(_0590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3413_ (.A(_2251_),
    .B(\ppwm_i.u_ppwm.global_counter[10] ),
    .C(_0590_),
    .Y(_0591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3414_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net784),
    .C1(_0591_),
    .B1(_2266_),
    .A1(\ppwm_i.u_ppwm.pwm_value[2] ),
    .Y(_0592_),
    .A2(_2265_));
 sg13g2_a221oi_1 _3415_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2250_),
    .C1(_0592_),
    .B1(\ppwm_i.u_ppwm.global_counter[12] ),
    .A1(_2249_),
    .Y(_0593_),
    .A2(\ppwm_i.u_ppwm.global_counter[13] ));
 sg13g2_a221oi_1 _3416_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.pwm_value[3] ),
    .C1(_0593_),
    .B1(_2264_),
    .A1(\ppwm_i.u_ppwm.pwm_value[4] ),
    .Y(_0594_),
    .A2(_2263_));
 sg13g2_a221oi_1 _3417_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2248_),
    .C1(_0594_),
    .B1(\ppwm_i.u_ppwm.global_counter[14] ),
    .A1(_2247_),
    .Y(_0595_),
    .A2(\ppwm_i.u_ppwm.global_counter[15] ));
 sg13g2_a221oi_1 _3418_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.pwm_value[5] ),
    .C1(_0595_),
    .B1(_2262_),
    .A1(\ppwm_i.u_ppwm.pwm_value[6] ),
    .Y(_0596_),
    .A2(_2261_));
 sg13g2_a221oi_1 _3419_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_2246_),
    .C1(_0596_),
    .B1(\ppwm_i.u_ppwm.global_counter[16] ),
    .A1(_2245_),
    .Y(_0597_),
    .A2(\ppwm_i.u_ppwm.global_counter[17] ));
 sg13g2_a221oi_1 _3420_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\ppwm_i.u_ppwm.pwm_value[7] ),
    .C1(_0597_),
    .B1(_2260_),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .Y(_0598_),
    .A2(_2259_));
 sg13g2_a21oi_1 _3421_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2244_),
    .A2(\ppwm_i.u_ppwm.global_counter[18] ),
    .Y(_0599_),
    .B1(_0598_));
 sg13g2_nor2_1 _3422_ (.A(_2243_),
    .B(\ppwm_i.u_ppwm.global_counter[19] ),
    .Y(_0600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3423_ (.B1(_0589_),
    .VDD(VPWR),
    .Y(_0601_),
    .VSS(VGND),
    .A1(_0599_),
    .A2(_0600_));
 sg13g2_nand3_1 _3424_ (.B(_0588_),
    .C(_0601_),
    .A(net610),
    .Y(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3425_ (.Y(_0603_),
    .A(_2419_),
    .B(_0602_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3426_ (.B1(_0532_),
    .VDD(VPWR),
    .Y(_0604_),
    .VSS(VGND),
    .A1(_0570_),
    .A2(_0603_));
 sg13g2_mux2_1 _3427_ (.A0(_0604_),
    .A1(net1162),
    .S(_0516_),
    .X(_0605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3428_ (.A(net821),
    .B(_0605_),
    .X(_0070_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _3429_ (.B(_2361_),
    .C(_2375_),
    .A(net419),
    .Y(_0606_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net582));
 sg13g2_o21ai_1 _3430_ (.B1(net813),
    .VDD(VPWR),
    .Y(_0607_),
    .VSS(VGND),
    .A1(net592),
    .A2(_0606_));
 sg13g2_a21oi_1 _3431_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2252_),
    .A2(_0606_),
    .Y(_0071_),
    .B1(_0607_));
 sg13g2_and2_1 _3432_ (.A(_2345_),
    .B(_2360_),
    .X(_0608_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3433_ (.A(net598),
    .B(net608),
    .Y(_0609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3434_ (.A(net608),
    .B_N(net611),
    .Y(_0610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3435_ (.B1(net579),
    .VDD(VPWR),
    .Y(_0611_),
    .VSS(VGND),
    .A1(_0609_),
    .A2(net589));
 sg13g2_nor2_1 _3436_ (.A(_2345_),
    .B(_2360_),
    .Y(_0612_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3437_ (.Y(_0613_),
    .B(_0612_),
    .A_N(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3438_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2255_),
    .Y(_0614_),
    .A2(_0613_),
    .A1(_0611_));
 sg13g2_a21o_1 _3439_ (.A2(_0613_),
    .A1(_0611_),
    .B1(_2255_),
    .X(_0615_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3440_ (.A(_2329_),
    .B(_2360_),
    .Y(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3441_ (.A(_2344_),
    .B(_0616_),
    .X(_0617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3442_ (.Y(_0618_),
    .A(_2344_),
    .B(_0616_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3443_ (.Y(_0619_),
    .A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3444_ (.Y(_0620_),
    .B(_0616_),
    .A_N(_2344_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3445_ (.Y(_0621_),
    .B(_2419_),
    .A_N(_0620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3446_ (.A(_2375_),
    .B(_0621_),
    .Y(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3447_ (.Y(_0623_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .B(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3448_ (.B1(_0623_),
    .VDD(VPWR),
    .Y(_0624_),
    .VSS(VGND),
    .A1(_2248_),
    .A2(net594));
 sg13g2_nand2_1 _3449_ (.Y(_0625_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .B(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3450_ (.B1(_0625_),
    .VDD(VPWR),
    .Y(_0626_),
    .VSS(VGND),
    .A1(_2249_),
    .A2(net595));
 sg13g2_mux2_1 _3451_ (.A0(_0626_),
    .A1(_0624_),
    .S(net609),
    .X(_0627_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3452_ (.A(net602),
    .B(_0621_),
    .Y(_0628_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3453_ (.A(net784),
    .B(net598),
    .Y(_0629_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3454_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2242_),
    .A2(net598),
    .Y(_0630_),
    .B1(_0629_));
 sg13g2_inv_1 _3455_ (.VDD(VPWR),
    .Y(_0631_),
    .A(_0630_),
    .VSS(VGND));
 sg13g2_nor2_1 _3456_ (.A(\ppwm_i.u_ppwm.pwm_value[2] ),
    .B(net595),
    .Y(_0632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3457_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0632_),
    .Y(_0633_),
    .A2(net595),
    .A1(_2241_));
 sg13g2_nand2_1 _3458_ (.Y(_0634_),
    .A(net611),
    .B(_0633_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3459_ (.B1(_0634_),
    .VDD(VPWR),
    .Y(_0635_),
    .VSS(VGND),
    .A1(net611),
    .A2(_0631_));
 sg13g2_a22oi_1 _3460_ (.Y(_0636_),
    .B1(net571),
    .B2(_0635_),
    .A2(_0627_),
    .A1(_0622_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3461_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0637_),
    .B(_0616_),
    .A(net579));
 sg13g2_nor2_1 _3462_ (.A(_2419_),
    .B(_0637_),
    .Y(_0638_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3463_ (.A(net594),
    .B_N(\ppwm_i.u_ppwm.global_counter[0] ),
    .Y(_0639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3464_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[10] ),
    .A2(net595),
    .Y(_0640_),
    .B1(_0639_));
 sg13g2_o21ai_1 _3465_ (.B1(net579),
    .VDD(VPWR),
    .Y(_0641_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .A2(net589));
 sg13g2_a21oi_1 _3466_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net589),
    .A2(_0640_),
    .Y(_0642_),
    .B1(_0641_));
 sg13g2_xnor2_1 _3467_ (.Y(_0643_),
    .A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3468_ (.A(_0618_),
    .B(_0643_),
    .Y(_0644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3469_ (.A(net573),
    .B(_0638_),
    .C(_0642_),
    .D(_0644_),
    .Y(_0645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3470_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0645_),
    .C1(net799),
    .B1(_0636_),
    .A1(_2251_),
    .Y(_0072_),
    .A2(net573));
 sg13g2_nand2_1 _3471_ (.Y(_0646_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3472_ (.B1(_0646_),
    .VDD(VPWR),
    .Y(_0647_),
    .VSS(VGND),
    .A1(_2247_),
    .A2(net596));
 sg13g2_mux2_1 _3473_ (.A0(_0624_),
    .A1(_0647_),
    .S(net609),
    .X(_0648_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3474_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0649_),
    .B(_0620_),
    .A(_2419_));
 sg13g2_nor2_1 _3475_ (.A(_2251_),
    .B(net598),
    .Y(_0650_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _3476_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_0650_),
    .Y(_0651_),
    .A2(net598),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ));
 sg13g2_nor3_1 _3477_ (.A(net584),
    .B(net574),
    .C(_0651_),
    .Y(_0652_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3478_ (.A(net609),
    .B_N(_0633_),
    .Y(_0653_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3479_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net609),
    .A2(_0626_),
    .Y(_0654_),
    .B1(_0653_));
 sg13g2_inv_1 _3480_ (.VDD(VPWR),
    .Y(_0655_),
    .A(_0654_),
    .VSS(VGND));
 sg13g2_a221oi_1 _3481_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net571),
    .C1(_0652_),
    .B1(_0655_),
    .A1(_0622_),
    .Y(_0656_),
    .A2(_0648_));
 sg13g2_nand2_1 _3482_ (.Y(_0657_),
    .A(net785),
    .B(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3483_ (.Y(_0658_),
    .A(net785),
    .B(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3484_ (.B1(net576),
    .VDD(VPWR),
    .Y(_0659_),
    .VSS(VGND),
    .A1(_0619_),
    .A2(_0658_));
 sg13g2_a21oi_1 _3485_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0619_),
    .A2(_0658_),
    .Y(_0660_),
    .B1(_0659_));
 sg13g2_nor2b_1 _3486_ (.A(net594),
    .B_N(\ppwm_i.u_ppwm.global_counter[1] ),
    .Y(_0661_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3487_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[11] ),
    .A2(net594),
    .Y(_0662_),
    .B1(_0661_));
 sg13g2_o21ai_1 _3488_ (.B1(net579),
    .VDD(VPWR),
    .Y(_0663_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .A2(net589));
 sg13g2_a21oi_1 _3489_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net589),
    .A2(_0662_),
    .Y(_0664_),
    .B1(_0663_));
 sg13g2_nor3_1 _3490_ (.A(_2381_),
    .B(_2388_),
    .C(_0637_),
    .Y(_0665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3491_ (.A(net573),
    .B(_0660_),
    .C(_0664_),
    .D(_0665_),
    .Y(_0666_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3492_ (.B1(net821),
    .VDD(VPWR),
    .Y(_0667_),
    .VSS(VGND),
    .A1(net784),
    .A2(_0614_));
 sg13g2_a21oi_1 _3493_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0656_),
    .A2(_0666_),
    .Y(_0073_),
    .B1(_0667_));
 sg13g2_xnor2_1 _3494_ (.Y(_0668_),
    .A(_2250_),
    .B(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3495_ (.B1(_0657_),
    .VDD(VPWR),
    .Y(_0669_),
    .VSS(VGND),
    .A1(_0619_),
    .A2(_0658_));
 sg13g2_nand2_1 _3496_ (.Y(_0670_),
    .A(_0668_),
    .B(_0669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3497_ (.A(net575),
    .B(_0670_),
    .X(_0671_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3498_ (.B1(_0671_),
    .VDD(VPWR),
    .Y(_0672_),
    .VSS(VGND),
    .A1(_0668_),
    .A2(_0669_));
 sg13g2_nand2_1 _3499_ (.Y(_0673_),
    .A(net611),
    .B(_0651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3500_ (.B1(_0673_),
    .VDD(VPWR),
    .Y(_0674_),
    .VSS(VGND),
    .A1(net584),
    .A2(_0630_));
 sg13g2_nor3_1 _3501_ (.A(net602),
    .B(net574),
    .C(_0674_),
    .Y(_0675_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3502_ (.Y(_0676_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3503_ (.B1(_0676_),
    .VDD(VPWR),
    .Y(_0677_),
    .VSS(VGND),
    .A1(_2246_),
    .A2(net597));
 sg13g2_mux2_1 _3504_ (.A0(_0647_),
    .A1(_0677_),
    .S(net610),
    .X(_0678_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3505_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0622_),
    .C1(_0675_),
    .B1(_0678_),
    .A1(_0627_),
    .Y(_0679_),
    .A2(net571));
 sg13g2_nor2_1 _3506_ (.A(net586),
    .B(_0637_),
    .Y(_0680_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3507_ (.A(_2272_),
    .B(net594),
    .Y(_0681_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3508_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[12] ),
    .A2(net594),
    .Y(_0682_),
    .B1(_0681_));
 sg13g2_o21ai_1 _3509_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0683_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .A2(net588));
 sg13g2_a21oi_1 _3510_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(_0682_),
    .Y(_0684_),
    .B1(_0683_));
 sg13g2_nor3_1 _3511_ (.A(net573),
    .B(_0680_),
    .C(_0684_),
    .Y(_0685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3512_ (.B(_0679_),
    .C(_0685_),
    .A(_0672_),
    .Y(_0686_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3513_ (.B1(_0686_),
    .VDD(VPWR),
    .Y(_0687_),
    .VSS(VGND),
    .A1(net1171),
    .A2(_0614_));
 sg13g2_nor2_1 _3514_ (.A(net798),
    .B(_0687_),
    .Y(_0074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3515_ (.B1(_0670_),
    .VDD(VPWR),
    .Y(_0688_),
    .VSS(VGND),
    .A1(_2250_),
    .A2(net586));
 sg13g2_nor2_1 _3516_ (.A(_2249_),
    .B(net586),
    .Y(_0689_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3517_ (.Y(_0690_),
    .A(_2249_),
    .B(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3518_ (.A(_0689_),
    .B_N(_0690_),
    .Y(_0691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3519_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0688_),
    .A2(_0691_),
    .Y(_0692_),
    .B1(_0618_));
 sg13g2_o21ai_1 _3520_ (.B1(_0692_),
    .VDD(VPWR),
    .Y(_0693_),
    .VSS(VGND),
    .A1(_0688_),
    .A2(_0691_));
 sg13g2_nand2_2 _3521_ (.Y(_0694_),
    .A(net602),
    .B(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3522_ (.VDD(VPWR),
    .Y(_0695_),
    .A(_0694_),
    .VSS(VGND));
 sg13g2_a22oi_1 _3523_ (.Y(_0696_),
    .B1(_0651_),
    .B2(net602),
    .A2(_0631_),
    .A1(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3524_ (.B1(_0696_),
    .VDD(VPWR),
    .Y(_0697_),
    .VSS(VGND),
    .A1(net584),
    .A2(_0633_));
 sg13g2_nor3_1 _3525_ (.A(net574),
    .B(_0695_),
    .C(_0697_),
    .Y(_0698_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3526_ (.Y(_0699_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .B(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3527_ (.B1(_0699_),
    .VDD(VPWR),
    .Y(_0700_),
    .VSS(VGND),
    .A1(_2245_),
    .A2(net597));
 sg13g2_mux2_1 _3528_ (.A0(_0677_),
    .A1(_0700_),
    .S(net610),
    .X(_0701_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3529_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0622_),
    .C1(_0698_),
    .B1(_0701_),
    .A1(net571),
    .Y(_0702_),
    .A2(_0648_));
 sg13g2_nand2_1 _3530_ (.Y(_0703_),
    .A(\ppwm_i.u_ppwm.global_counter[13] ),
    .B(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3531_ (.B1(_0703_),
    .VDD(VPWR),
    .Y(_0704_),
    .VSS(VGND),
    .A1(_2271_),
    .A2(net593));
 sg13g2_mux2_1 _3532_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .A1(_0704_),
    .S(net588),
    .X(_0705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3533_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_0705_),
    .Y(_0706_),
    .B1(net572));
 sg13g2_and2_1 _3534_ (.A(_0702_),
    .B(_0706_),
    .X(_0707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3535_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0707_),
    .C1(net798),
    .B1(_0693_),
    .A1(_2249_),
    .Y(_0075_),
    .A2(net572));
 sg13g2_nor2_1 _3536_ (.A(_2248_),
    .B(net586),
    .Y(_0708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3537_ (.Y(_0709_),
    .A(_2248_),
    .B(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3538_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0688_),
    .A2(_0690_),
    .Y(_0710_),
    .B1(_0689_));
 sg13g2_nor2b_1 _3539_ (.A(_0709_),
    .B_N(_0710_),
    .Y(_0711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3540_ (.A(_0710_),
    .B_N(_0709_),
    .Y(_0712_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3541_ (.A(_0618_),
    .B(_0711_),
    .C(_0712_),
    .Y(_0713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _3542_ (.Y(_0714_),
    .A(net584),
    .B(_0694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3543_ (.A(_0635_),
    .B(_0714_),
    .Y(_0715_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3544_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0651_),
    .A2(_0695_),
    .Y(_0716_),
    .B1(net574));
 sg13g2_o21ai_1 _3545_ (.B1(_0716_),
    .VDD(VPWR),
    .Y(_0717_),
    .VSS(VGND),
    .A1(net584),
    .A2(_0626_));
 sg13g2_nand2_1 _3546_ (.Y(_0718_),
    .A(net782),
    .B(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3547_ (.B1(_0718_),
    .VDD(VPWR),
    .Y(_0719_),
    .VSS(VGND),
    .A1(_2244_),
    .A2(net599));
 sg13g2_mux2_1 _3548_ (.A0(_0700_),
    .A1(_0719_),
    .S(net609),
    .X(_0720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3549_ (.Y(_0721_),
    .B1(_0720_),
    .B2(_0622_),
    .A2(_0678_),
    .A1(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3550_ (.B1(_0721_),
    .VDD(VPWR),
    .Y(_0722_),
    .VSS(VGND),
    .A1(_0715_),
    .A2(_0717_));
 sg13g2_nor2_1 _3551_ (.A(_2270_),
    .B(net593),
    .Y(_0723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3552_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net974),
    .A2(net593),
    .Y(_0724_),
    .B1(_0723_));
 sg13g2_o21ai_1 _3553_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0725_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .A2(net588));
 sg13g2_a21oi_1 _3554_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(_0724_),
    .Y(_0726_),
    .B1(_0725_));
 sg13g2_nor4_1 _3555_ (.A(net572),
    .B(_0713_),
    .C(_0722_),
    .D(_0726_),
    .Y(_0727_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3556_ (.B1(net822),
    .VDD(VPWR),
    .Y(_0728_),
    .VSS(VGND),
    .A1(net1181),
    .A2(_0614_));
 sg13g2_nor2_1 _3557_ (.A(_0727_),
    .B(_0728_),
    .Y(_0076_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3558_ (.Y(_0729_),
    .A(_2247_),
    .B(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _3559_ (.A(_0708_),
    .B(_0712_),
    .C(_0729_),
    .X(_0730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3560_ (.B1(_0729_),
    .VDD(VPWR),
    .Y(_0731_),
    .VSS(VGND),
    .A1(_0708_),
    .A2(_0712_));
 sg13g2_nand3_1 _3561_ (.B(_0730_),
    .C(_0731_),
    .A(net575),
    .Y(_0732_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3562_ (.A(_0655_),
    .B(_0714_),
    .Y(_0733_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3563_ (.A(_0630_),
    .B(_0694_),
    .Y(_0734_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3564_ (.A(net584),
    .B(_0624_),
    .Y(_0735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3565_ (.A(net574),
    .B(_0733_),
    .C(_0734_),
    .D(_0735_),
    .Y(_0736_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3566_ (.A(net609),
    .B(_0719_),
    .Y(_0737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3567_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .A2(net596),
    .Y(_0738_),
    .B1(_0548_));
 sg13g2_a21oi_1 _3568_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net610),
    .A2(_0738_),
    .Y(_0739_),
    .B1(_0737_));
 sg13g2_a221oi_1 _3569_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0622_),
    .C1(_0736_),
    .B1(_0739_),
    .A1(net571),
    .Y(_0740_),
    .A2(_0701_));
 sg13g2_nor2_1 _3570_ (.A(\ppwm_i.u_ppwm.global_counter[5] ),
    .B(net593),
    .Y(_0741_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3571_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2262_),
    .A2(net593),
    .Y(_0742_),
    .B1(_0741_));
 sg13g2_mux2_1 _3572_ (.A0(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .A1(_0742_),
    .S(net588),
    .X(_0743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3573_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net578),
    .A2(_0743_),
    .Y(_0744_),
    .B1(net572));
 sg13g2_and2_1 _3574_ (.A(_0740_),
    .B(_0744_),
    .X(_0745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3575_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0745_),
    .C1(net799),
    .B1(_0732_),
    .A1(_2247_),
    .Y(_0077_),
    .A2(net572));
 sg13g2_xnor2_1 _3576_ (.Y(_0746_),
    .A(_2246_),
    .B(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3577_ (.B1(net600),
    .VDD(VPWR),
    .Y(_0747_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[5] ),
    .A2(\ppwm_i.u_ppwm.pwm_value[4] ));
 sg13g2_nand2_1 _3578_ (.Y(_0748_),
    .A(_0712_),
    .B(_0729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3579_ (.Y(_0749_),
    .A(_0747_),
    .B(_0748_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3580_ (.A(_0746_),
    .B(_0749_),
    .X(_0750_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3581_ (.A(_0618_),
    .B(_0750_),
    .Y(_0751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3582_ (.B1(_0751_),
    .VDD(VPWR),
    .Y(_0752_),
    .VSS(VGND),
    .A1(_0746_),
    .A2(_0749_));
 sg13g2_nor2_1 _3583_ (.A(_0633_),
    .B(_0694_),
    .Y(_0753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3584_ (.A(net584),
    .B(_0647_),
    .Y(_0754_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _3585_ (.A(net574),
    .B(_0753_),
    .C(_0754_),
    .Y(_0755_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3586_ (.B1(_0755_),
    .VDD(VPWR),
    .Y(_0756_),
    .VSS(VGND),
    .A1(_0627_),
    .A2(_0714_));
 sg13g2_nor2_1 _3587_ (.A(net609),
    .B(_0738_),
    .Y(_0757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3588_ (.Y(_0758_),
    .B1(_0757_),
    .B2(_0622_),
    .A2(_0720_),
    .A1(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3589_ (.Y(_0759_),
    .A(_0756_),
    .B(_0758_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3590_ (.A(_2269_),
    .B(net592),
    .Y(_0760_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3591_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[16] ),
    .A2(net592),
    .Y(_0761_),
    .B1(_0760_));
 sg13g2_o21ai_1 _3592_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0762_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .A2(net588));
 sg13g2_a21oi_1 _3593_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net588),
    .A2(_0761_),
    .Y(_0763_),
    .B1(_0762_));
 sg13g2_nor3_1 _3594_ (.A(net572),
    .B(_0759_),
    .C(_0763_),
    .Y(_0764_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3595_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0764_),
    .C1(net798),
    .B1(_0752_),
    .A1(_2246_),
    .Y(_0078_),
    .A2(net572));
 sg13g2_xnor2_1 _3596_ (.Y(_0765_),
    .A(_2245_),
    .B(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3597_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1187),
    .A2(net601),
    .Y(_0766_),
    .B1(_0750_));
 sg13g2_nand2b_1 _3598_ (.Y(_0767_),
    .B(_0766_),
    .A_N(_0765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3599_ (.Y(_0768_),
    .B(_0765_),
    .A_N(_0766_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3600_ (.B(_0767_),
    .C(_0768_),
    .A(net575),
    .Y(_0769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3601_ (.A(net584),
    .B(_0677_),
    .Y(_0770_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3602_ (.A(_0626_),
    .B(_0694_),
    .Y(_0771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3603_ (.A(_0648_),
    .B(_0714_),
    .Y(_0772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3604_ (.A(_0649_),
    .B(_0770_),
    .C(_0771_),
    .D(_0772_),
    .Y(_0773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3605_ (.A2(_0739_),
    .A1(net571),
    .B1(_0773_),
    .X(_0774_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3606_ (.A(_2268_),
    .B(net592),
    .Y(_0775_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3607_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.global_counter[17] ),
    .A2(net591),
    .Y(_0776_),
    .B1(_0775_));
 sg13g2_o21ai_1 _3608_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0777_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .A2(net590));
 sg13g2_a21oi_1 _3609_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net590),
    .A2(_0776_),
    .Y(_0778_),
    .B1(_0777_));
 sg13g2_nor3_1 _3610_ (.A(net572),
    .B(_0774_),
    .C(_0778_),
    .Y(_0779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3611_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0779_),
    .C1(net798),
    .B1(_0769_),
    .A1(_2245_),
    .Y(_0079_),
    .A2(net573));
 sg13g2_nand4_1 _3612_ (.B(_0729_),
    .C(_0746_),
    .A(_0712_),
    .Y(_0780_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0765_));
 sg13g2_o21ai_1 _3613_ (.B1(net601),
    .VDD(VPWR),
    .Y(_0781_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[7] ),
    .A2(\ppwm_i.u_ppwm.pwm_value[6] ));
 sg13g2_and3_2 _3614_ (.X(_0782_),
    .A(_0747_),
    .B(_0780_),
    .C(_0781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3615_ (.Y(_0783_),
    .A(_2244_),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3616_ (.Y(_0784_),
    .B(_0782_),
    .A_N(_0783_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _3617_ (.A(_0782_),
    .B_N(_0783_),
    .Y(_0785_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _3618_ (.B(net576),
    .C(_0784_),
    .Y(_0786_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0785_));
 sg13g2_nor2_1 _3619_ (.A(net585),
    .B(_0700_),
    .Y(_0787_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3620_ (.A(_0624_),
    .B(_0694_),
    .Y(_0788_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3621_ (.A(_0678_),
    .B(_0714_),
    .Y(_0789_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3622_ (.A(net574),
    .B(_0787_),
    .C(_0788_),
    .D(_0789_),
    .Y(_0790_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3623_ (.A2(_0757_),
    .A1(_0628_),
    .B1(_0790_),
    .X(_0791_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3624_ (.Y(_0792_),
    .A(\ppwm_i.u_ppwm.global_counter[18] ),
    .B(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3625_ (.B1(_0792_),
    .VDD(VPWR),
    .Y(_0793_),
    .VSS(VGND),
    .A1(_2267_),
    .A2(net591));
 sg13g2_inv_1 _3626_ (.VDD(VPWR),
    .Y(_0794_),
    .A(_0793_),
    .VSS(VGND));
 sg13g2_o21ai_1 _3627_ (.B1(net580),
    .VDD(VPWR),
    .Y(_0795_),
    .VSS(VGND),
    .A1(net783),
    .A2(net589));
 sg13g2_a21oi_1 _3628_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net589),
    .A2(_0794_),
    .Y(_0796_),
    .B1(_0795_));
 sg13g2_nor3_1 _3629_ (.A(net573),
    .B(_0791_),
    .C(_0796_),
    .Y(_0797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3630_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0797_),
    .C1(net799),
    .B1(_0786_),
    .A1(_2244_),
    .Y(_0080_),
    .A2(net573));
 sg13g2_a21oi_1 _3631_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .A2(net603),
    .Y(_0798_),
    .B1(_0785_));
 sg13g2_xnor2_1 _3632_ (.Y(_0799_),
    .A(\ppwm_i.u_ppwm.pwm_value[9] ),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3633_ (.B1(net576),
    .VDD(VPWR),
    .Y(_0800_),
    .VSS(VGND),
    .A1(_0798_),
    .A2(_0799_));
 sg13g2_a21oi_1 _3634_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0798_),
    .A2(_0799_),
    .Y(_0801_),
    .B1(_0800_));
 sg13g2_nor2_1 _3635_ (.A(net585),
    .B(_0719_),
    .Y(_0802_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3636_ (.A(_0647_),
    .B(_0694_),
    .Y(_0803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3637_ (.A(_0701_),
    .B(_0714_),
    .Y(_0804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _3638_ (.A(net574),
    .B(_0802_),
    .C(_0803_),
    .D(_0804_),
    .Y(_0805_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3639_ (.B1(_0586_),
    .VDD(VPWR),
    .Y(_0806_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.global_counter[9] ),
    .A2(net592));
 sg13g2_o21ai_1 _3640_ (.B1(net579),
    .VDD(VPWR),
    .Y(_0807_),
    .VSS(VGND),
    .A1(net1160),
    .A2(net589));
 sg13g2_a21oi_1 _3641_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net590),
    .A2(_0806_),
    .Y(_0808_),
    .B1(_0807_));
 sg13g2_nor4_1 _3642_ (.A(_0615_),
    .B(_0801_),
    .C(_0805_),
    .D(_0808_),
    .Y(_0809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3643_ (.B1(net821),
    .VDD(VPWR),
    .Y(_0810_),
    .VSS(VGND),
    .A1(net1167),
    .A2(_0614_));
 sg13g2_nor2_1 _3644_ (.A(_0809_),
    .B(_0810_),
    .Y(_0081_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3645_ (.A(net612),
    .B(_0609_),
    .Y(_0811_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _3646_ (.Y(_0812_),
    .B1(_0811_),
    .B2(net579),
    .A2(_0612_),
    .A1(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3647_ (.A(_2255_),
    .B(_0812_),
    .Y(_0813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _3648_ (.Y(_0814_),
    .B(net419),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_0812_));
 sg13g2_nand2_1 _3649_ (.Y(_0815_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .B(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3650_ (.A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .B(net582),
    .Y(_0816_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3651_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net582),
    .A2(_0640_),
    .Y(_0817_),
    .B1(_0816_));
 sg13g2_xor2_1 _3652_ (.B(net608),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .X(_0818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3653_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net576),
    .C1(_0638_),
    .B1(_0818_),
    .A1(net579),
    .Y(_0819_),
    .A2(_0817_));
 sg13g2_nand3_1 _3654_ (.B(_0813_),
    .C(_0819_),
    .A(_0636_),
    .Y(_0820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3655_ (.B1(_0820_),
    .VDD(VPWR),
    .Y(_0821_),
    .VSS(VGND),
    .A1(net1173),
    .A2(_0813_));
 sg13g2_nor2_1 _3656_ (.A(net799),
    .B(_0821_),
    .Y(_0082_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3657_ (.Y(_0822_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .B(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3658_ (.Y(_0823_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .B(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _3659_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0824_),
    .B(_0823_),
    .A(_0815_));
 sg13g2_a21oi_1 _3660_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0815_),
    .A2(_0823_),
    .Y(_0825_),
    .B1(_0618_));
 sg13g2_and2_1 _3661_ (.A(_0824_),
    .B(_0825_),
    .X(_0826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3662_ (.B1(net579),
    .VDD(VPWR),
    .Y(_0827_),
    .VSS(VGND),
    .A1(net785),
    .A2(net582));
 sg13g2_a21oi_1 _3663_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net582),
    .A2(_0662_),
    .Y(_0828_),
    .B1(_0827_));
 sg13g2_nor4_1 _3664_ (.A(_0665_),
    .B(net570),
    .C(_0826_),
    .D(_0828_),
    .Y(_0829_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3665_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0656_),
    .C1(net799),
    .B1(_0829_),
    .A1(_2242_),
    .Y(_0083_),
    .A2(net570));
 sg13g2_xnor2_1 _3666_ (.Y(_0830_),
    .A(_2241_),
    .B(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3667_ (.VDD(VPWR),
    .Y(_0831_),
    .A(_0830_),
    .VSS(VGND));
 sg13g2_a21o_1 _3668_ (.A2(_0824_),
    .A1(_0822_),
    .B1(_0831_),
    .X(_0832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3669_ (.B(_0824_),
    .C(_0831_),
    .A(_0822_),
    .Y(_0833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _3670_ (.X(_0834_),
    .A(net576),
    .B(_0832_),
    .C(_0833_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3671_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0835_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[2] ),
    .A2(net582));
 sg13g2_a21oi_1 _3672_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net582),
    .A2(_0682_),
    .Y(_0836_),
    .B1(_0835_));
 sg13g2_nor4_1 _3673_ (.A(_0680_),
    .B(net570),
    .C(_0834_),
    .D(_0836_),
    .Y(_0837_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3674_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0679_),
    .C1(net798),
    .B1(_0837_),
    .A1(_2241_),
    .Y(_0084_),
    .A2(net570));
 sg13g2_o21ai_1 _3675_ (.B1(_0832_),
    .VDD(VPWR),
    .Y(_0838_),
    .VSS(VGND),
    .A1(_2241_),
    .A2(net586));
 sg13g2_nor2_1 _3676_ (.A(_2240_),
    .B(net586),
    .Y(_0839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3677_ (.Y(_0840_),
    .A(_2240_),
    .B(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3678_ (.Y(_0841_),
    .B(_0840_),
    .A_N(_0839_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3679_ (.Y(_0842_),
    .A(_0838_),
    .B(_0841_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _3680_ (.A0(\ppwm_i.u_ppwm.pwm_value[3] ),
    .A1(_0704_),
    .S(net581),
    .X(_0843_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3681_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net577),
    .A2(_0843_),
    .Y(_0844_),
    .B1(net569));
 sg13g2_nand2_1 _3682_ (.Y(_0845_),
    .A(_0702_),
    .B(_0844_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3683_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net575),
    .A2(_0842_),
    .Y(_0846_),
    .B1(_0845_));
 sg13g2_o21ai_1 _3684_ (.B1(net822),
    .VDD(VPWR),
    .Y(_0847_),
    .VSS(VGND),
    .A1(net1151),
    .A2(_0813_));
 sg13g2_nor2_1 _3685_ (.A(_0846_),
    .B(_0847_),
    .Y(_0085_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3686_ (.Y(_0848_),
    .A(_2239_),
    .B(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3687_ (.A2(_0840_),
    .A1(_0838_),
    .B1(_0839_),
    .X(_0849_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3688_ (.A(_0848_),
    .B(_0849_),
    .X(_0850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3689_ (.A(_0618_),
    .B(_0850_),
    .Y(_0851_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3690_ (.B1(_0851_),
    .VDD(VPWR),
    .Y(_0852_),
    .VSS(VGND),
    .A1(_0848_),
    .A2(_0849_));
 sg13g2_o21ai_1 _3691_ (.B1(net577),
    .VDD(VPWR),
    .Y(_0853_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[4] ),
    .A2(net581));
 sg13g2_a21oi_1 _3692_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net581),
    .A2(_0724_),
    .Y(_0854_),
    .B1(_0853_));
 sg13g2_nor3_1 _3693_ (.A(_0722_),
    .B(net569),
    .C(_0854_),
    .Y(_0855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3694_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0855_),
    .C1(net795),
    .B1(_0852_),
    .A1(_2239_),
    .Y(_0086_),
    .A2(net569));
 sg13g2_xnor2_1 _3695_ (.Y(_0856_),
    .A(_2238_),
    .B(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _3696_ (.VDD(VPWR),
    .Y(_0857_),
    .A(_0856_),
    .VSS(VGND));
 sg13g2_a21oi_1 _3697_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .A2(net600),
    .Y(_0858_),
    .B1(_0850_));
 sg13g2_a21oi_1 _3698_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_0857_),
    .A2(_0858_),
    .Y(_0859_),
    .B1(_0618_));
 sg13g2_o21ai_1 _3699_ (.B1(_0859_),
    .VDD(VPWR),
    .Y(_0860_),
    .VSS(VGND),
    .A1(_0857_),
    .A2(_0858_));
 sg13g2_mux2_1 _3700_ (.A0(\ppwm_i.u_ppwm.pwm_value[5] ),
    .A1(_0742_),
    .S(net581),
    .X(_0861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3701_ (.Y(_0862_),
    .A(_0740_),
    .B(_0813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3702_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net578),
    .A2(_0861_),
    .Y(_0863_),
    .B1(_0862_));
 sg13g2_a221oi_1 _3703_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0863_),
    .C1(net795),
    .B1(_0860_),
    .A1(_2238_),
    .Y(_0087_),
    .A2(net569));
 sg13g2_xnor2_1 _3704_ (.Y(_0864_),
    .A(_2237_),
    .B(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3705_ (.B1(net600),
    .VDD(VPWR),
    .Y(_0865_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .A2(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ));
 sg13g2_nand2_1 _3706_ (.Y(_0866_),
    .A(_0850_),
    .B(_0856_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3707_ (.Y(_0867_),
    .A(_0865_),
    .B(_0866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3708_ (.A(_0864_),
    .B(_0867_),
    .X(_0868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3709_ (.B1(net575),
    .VDD(VPWR),
    .Y(_0869_),
    .VSS(VGND),
    .A1(_0864_),
    .A2(_0867_));
 sg13g2_or2_1 _3710_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_0870_),
    .B(_0869_),
    .A(_0868_));
 sg13g2_o21ai_1 _3711_ (.B1(net578),
    .VDD(VPWR),
    .Y(_0871_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[6] ),
    .A2(net581));
 sg13g2_a21oi_1 _3712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net581),
    .A2(_0761_),
    .Y(_0872_),
    .B1(_0871_));
 sg13g2_nor3_1 _3713_ (.A(_0759_),
    .B(net569),
    .C(_0872_),
    .Y(_0873_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3714_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0873_),
    .C1(net798),
    .B1(_0870_),
    .A1(_2237_),
    .Y(_0088_),
    .A2(net569));
 sg13g2_xnor2_1 _3715_ (.Y(_0874_),
    .A(_2236_),
    .B(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .A2(net601),
    .Y(_0875_),
    .B1(_0868_));
 sg13g2_nand2b_1 _3717_ (.Y(_0876_),
    .B(_0875_),
    .A_N(_0874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _3718_ (.Y(_0877_),
    .B(_0874_),
    .A_N(_0875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3719_ (.B(_0876_),
    .C(_0877_),
    .A(net575),
    .Y(_0878_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3720_ (.B1(net578),
    .VDD(VPWR),
    .Y(_0879_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[7] ),
    .A2(net583));
 sg13g2_a21oi_1 _3721_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net581),
    .A2(_0776_),
    .Y(_0880_),
    .B1(_0879_));
 sg13g2_nor3_1 _3722_ (.A(_0774_),
    .B(net569),
    .C(_0880_),
    .Y(_0881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3723_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0881_),
    .C1(net798),
    .B1(_0878_),
    .A1(_2236_),
    .Y(_0089_),
    .A2(net569));
 sg13g2_nand4_1 _3724_ (.B(_0856_),
    .C(_0864_),
    .A(_0850_),
    .Y(_0882_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_0874_));
 sg13g2_o21ai_1 _3725_ (.B1(net601),
    .VDD(VPWR),
    .Y(_0883_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .A2(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ));
 sg13g2_nand3_1 _3726_ (.B(_0882_),
    .C(_0883_),
    .A(_0865_),
    .Y(_0884_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3727_ (.Y(_0885_),
    .A(net783),
    .B(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _3728_ (.B(net602),
    .A(net783),
    .X(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3729_ (.Y(_0887_),
    .A(_0884_),
    .B(_0886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3730_ (.B1(net575),
    .VDD(VPWR),
    .Y(_0888_),
    .VSS(VGND),
    .A1(_0884_),
    .A2(_0886_));
 sg13g2_nor2b_1 _3731_ (.A(_0888_),
    .B_N(_0887_),
    .Y(_0889_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3732_ (.B1(net580),
    .VDD(VPWR),
    .Y(_0890_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[8] ),
    .A2(net583));
 sg13g2_a21oi_1 _3733_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net582),
    .A2(_0794_),
    .Y(_0891_),
    .B1(_0890_));
 sg13g2_nor4_1 _3734_ (.A(_0791_),
    .B(net570),
    .C(_0889_),
    .D(_0891_),
    .Y(_0892_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3735_ (.B1(net822),
    .VDD(VPWR),
    .Y(_0893_),
    .VSS(VGND),
    .A1(net783),
    .A2(_0813_));
 sg13g2_nor2_1 _3736_ (.A(_0892_),
    .B(_0893_),
    .Y(_0090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _3737_ (.Y(_0894_),
    .A(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .B(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3738_ (.B(_0887_),
    .C(_0894_),
    .A(_0885_),
    .Y(_0895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _3739_ (.A2(_0887_),
    .A1(_0885_),
    .B1(_0894_),
    .X(_0896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3740_ (.B(_0895_),
    .C(_0896_),
    .A(net575),
    .Y(_0897_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3741_ (.B1(net580),
    .VDD(VPWR),
    .Y(_0898_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.pwm_value[9] ),
    .A2(net583));
 sg13g2_a21oi_1 _3742_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net583),
    .A2(_0806_),
    .Y(_0899_),
    .B1(_0898_));
 sg13g2_nor3_1 _3743_ (.A(_0805_),
    .B(net570),
    .C(_0899_),
    .Y(_0900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _3744_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_0900_),
    .C1(net798),
    .B1(_0897_),
    .A1(_2235_),
    .Y(_0091_),
    .A2(net570));
 sg13g2_nand2_1 _3745_ (.Y(_0901_),
    .A(net459),
    .B(net1015),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _3746_ (.B(\falu_i.falutop.i2c_inst.state[0] ),
    .C(net804),
    .A(net459),
    .Y(_0902_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3747_ (.A(\falu_i.falutop.i2c_inst.data_in[16] ),
    .B(net686),
    .Y(_0903_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3748_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2291_),
    .A2(net685),
    .Y(_0092_),
    .B1(_0903_));
 sg13g2_mux2_1 _3749_ (.A0(net912),
    .A1(\falu_i.falutop.i2c_inst.op[1] ),
    .S(net686),
    .X(_0093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _3750_ (.A(\falu_i.falutop.i2c_inst.data_in[18] ),
    .B(net686),
    .Y(_0904_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3751_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2293_),
    .A2(net686),
    .Y(_0094_),
    .B1(_0904_));
 sg13g2_nor2_1 _3752_ (.A(\falu_i.falutop.i2c_inst.data_in[19] ),
    .B(net686),
    .Y(_0905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3753_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2292_),
    .A2(net686),
    .Y(_0095_),
    .B1(_0905_));
 sg13g2_and2_1 _3754_ (.A(net807),
    .B(net5),
    .X(_0096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3755_ (.A(net807),
    .B(net374),
    .X(_0097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3756_ (.A(net807),
    .B(net375),
    .X(_0098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3757_ (.A(net807),
    .B(net4),
    .X(_0099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _3758_ (.A(\ppwm_i.u_ppwm.u_mem.clk_prog_sync3 ),
    .B_N(net375),
    .Y(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3759_ (.A(net883),
    .B(_0906_),
    .X(_0907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3760_ (.Y(_0908_),
    .A(\ppwm_i.u_ppwm.u_mem.programming ),
    .B(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3761_ (.B1(net836),
    .VDD(VPWR),
    .Y(_0909_),
    .VSS(VGND),
    .A1(net868),
    .A2(net662));
 sg13g2_a21oi_1 _3762_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2234_),
    .A2(net662),
    .Y(_0100_),
    .B1(_0909_));
 sg13g2_o21ai_1 _3763_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0910_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[2] ),
    .A2(net644));
 sg13g2_a21oi_1 _3764_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2234_),
    .A2(net644),
    .Y(_0101_),
    .B1(_0910_));
 sg13g2_o21ai_1 _3765_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0911_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[2] ),
    .A2(net661));
 sg13g2_a21oi_1 _3766_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2233_),
    .A2(net661),
    .Y(_0102_),
    .B1(_0911_));
 sg13g2_o21ai_1 _3767_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0912_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[3] ),
    .A2(net659));
 sg13g2_a21oi_1 _3768_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2232_),
    .A2(net659),
    .Y(_0103_),
    .B1(_0912_));
 sg13g2_o21ai_1 _3769_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0913_),
    .VSS(VGND),
    .A1(net847),
    .A2(net642));
 sg13g2_a21oi_1 _3770_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2232_),
    .A2(net641),
    .Y(_0104_),
    .B1(_0913_));
 sg13g2_o21ai_1 _3771_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0914_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .A2(net655));
 sg13g2_a21oi_1 _3772_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2231_),
    .A2(net654),
    .Y(_0105_),
    .B1(_0914_));
 sg13g2_o21ai_1 _3773_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0915_),
    .VSS(VGND),
    .A1(net483),
    .A2(net654));
 sg13g2_a21oi_1 _3774_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2230_),
    .A2(net654),
    .Y(_0106_),
    .B1(_0915_));
 sg13g2_o21ai_1 _3775_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0916_),
    .VSS(VGND),
    .A1(net451),
    .A2(net662));
 sg13g2_a21oi_1 _3776_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2229_),
    .A2(net662),
    .Y(_0107_),
    .B1(_0916_));
 sg13g2_o21ai_1 _3777_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0917_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .A2(net644));
 sg13g2_a21oi_1 _3778_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2229_),
    .A2(net644),
    .Y(_0108_),
    .B1(_0917_));
 sg13g2_o21ai_1 _3779_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0918_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .A2(net662));
 sg13g2_a21oi_1 _3780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2228_),
    .A2(net662),
    .Y(_0109_),
    .B1(_0918_));
 sg13g2_o21ai_1 _3781_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0919_),
    .VSS(VGND),
    .A1(net504),
    .A2(net660));
 sg13g2_a21oi_1 _3782_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2227_),
    .A2(net660),
    .Y(_0110_),
    .B1(_0919_));
 sg13g2_o21ai_1 _3783_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0920_),
    .VSS(VGND),
    .A1(net888),
    .A2(net655));
 sg13g2_a21oi_1 _3784_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2226_),
    .A2(net655),
    .Y(_0111_),
    .B1(_0920_));
 sg13g2_o21ai_1 _3785_ (.B1(net832),
    .VDD(VPWR),
    .Y(_0921_),
    .VSS(VGND),
    .A1(net933),
    .A2(net641));
 sg13g2_a21oi_1 _3786_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2226_),
    .A2(net641),
    .Y(_0112_),
    .B1(_0921_));
 sg13g2_o21ai_1 _3787_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0922_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .A2(net653));
 sg13g2_a21oi_1 _3788_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2225_),
    .A2(net653),
    .Y(_0113_),
    .B1(_0922_));
 sg13g2_o21ai_1 _3789_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0923_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[14] ),
    .A2(net661));
 sg13g2_a21oi_1 _3790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2224_),
    .A2(net661),
    .Y(_0114_),
    .B1(_0923_));
 sg13g2_o21ai_1 _3791_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0924_),
    .VSS(VGND),
    .A1(net515),
    .A2(net644));
 sg13g2_a21oi_1 _3792_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2224_),
    .A2(net644),
    .Y(_0115_),
    .B1(_0924_));
 sg13g2_o21ai_1 _3793_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0925_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .A2(net659));
 sg13g2_a21oi_1 _3794_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2223_),
    .A2(net659),
    .Y(_0116_),
    .B1(_0925_));
 sg13g2_o21ai_1 _3795_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0926_),
    .VSS(VGND),
    .A1(net447),
    .A2(net659));
 sg13g2_a21oi_1 _3796_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2222_),
    .A2(net659),
    .Y(_0117_),
    .B1(_0926_));
 sg13g2_o21ai_1 _3797_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0927_),
    .VSS(VGND),
    .A1(net898),
    .A2(net653));
 sg13g2_a21oi_1 _3798_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2221_),
    .A2(net653),
    .Y(_0118_),
    .B1(_0927_));
 sg13g2_o21ai_1 _3799_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0928_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .A2(net641));
 sg13g2_a21oi_1 _3800_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2221_),
    .A2(net641),
    .Y(_0119_),
    .B1(_0928_));
 sg13g2_o21ai_1 _3801_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0929_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .A2(net653));
 sg13g2_a21oi_1 _3802_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2220_),
    .A2(net653),
    .Y(_0120_),
    .B1(_0929_));
 sg13g2_o21ai_1 _3803_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0930_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[21] ),
    .A2(net661));
 sg13g2_a21oi_1 _3804_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2219_),
    .A2(net661),
    .Y(_0121_),
    .B1(_0930_));
 sg13g2_o21ai_1 _3805_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0931_),
    .VSS(VGND),
    .A1(net844),
    .A2(net644));
 sg13g2_a21oi_1 _3806_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2219_),
    .A2(net644),
    .Y(_0122_),
    .B1(_0931_));
 sg13g2_o21ai_1 _3807_ (.B1(net828),
    .VDD(VPWR),
    .Y(_0932_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .A2(net661));
 sg13g2_a21oi_1 _3808_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2218_),
    .A2(net661),
    .Y(_0123_),
    .B1(_0932_));
 sg13g2_o21ai_1 _3809_ (.B1(net827),
    .VDD(VPWR),
    .Y(_0933_),
    .VSS(VGND),
    .A1(net402),
    .A2(net659));
 sg13g2_a21oi_1 _3810_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2217_),
    .A2(net659),
    .Y(_0124_),
    .B1(_0933_));
 sg13g2_o21ai_1 _3811_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0934_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[25] ),
    .A2(net653));
 sg13g2_a21oi_1 _3812_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2216_),
    .A2(net655),
    .Y(_0125_),
    .B1(_0934_));
 sg13g2_o21ai_1 _3813_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0935_),
    .VSS(VGND),
    .A1(net963),
    .A2(net641));
 sg13g2_a21oi_1 _3814_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2216_),
    .A2(net641),
    .Y(_0126_),
    .B1(_0935_));
 sg13g2_o21ai_1 _3815_ (.B1(net824),
    .VDD(VPWR),
    .Y(_0936_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .A2(net654));
 sg13g2_a21oi_1 _3816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2215_),
    .A2(net654),
    .Y(_0127_),
    .B1(_0936_));
 sg13g2_o21ai_1 _3817_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0937_),
    .VSS(VGND),
    .A1(net959),
    .A2(net660));
 sg13g2_a21oi_1 _3818_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2214_),
    .A2(net660),
    .Y(_0128_),
    .B1(_0937_));
 sg13g2_o21ai_1 _3819_ (.B1(net831),
    .VDD(VPWR),
    .Y(_0938_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .A2(net643));
 sg13g2_a21oi_1 _3820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2214_),
    .A2(net643),
    .Y(_0129_),
    .B1(_0938_));
 sg13g2_o21ai_1 _3821_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0939_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .A2(net664));
 sg13g2_a21oi_1 _3822_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2213_),
    .A2(net664),
    .Y(_0130_),
    .B1(_0939_));
 sg13g2_o21ai_1 _3823_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0940_),
    .VSS(VGND),
    .A1(net516),
    .A2(net656));
 sg13g2_a21oi_1 _3824_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2212_),
    .A2(net657),
    .Y(_0131_),
    .B1(_0940_));
 sg13g2_o21ai_1 _3825_ (.B1(net826),
    .VDD(VPWR),
    .Y(_0941_),
    .VSS(VGND),
    .A1(net534),
    .A2(net658));
 sg13g2_a21oi_1 _3826_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2211_),
    .A2(net658),
    .Y(_0132_),
    .B1(_0941_));
 sg13g2_o21ai_1 _3827_ (.B1(net826),
    .VDD(VPWR),
    .Y(_0942_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .A2(net642));
 sg13g2_a21oi_1 _3828_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2211_),
    .A2(net642),
    .Y(_0133_),
    .B1(_0942_));
 sg13g2_o21ai_1 _3829_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0943_),
    .VSS(VGND),
    .A1(net897),
    .A2(net656));
 sg13g2_a21oi_1 _3830_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2210_),
    .A2(net656),
    .Y(_0134_),
    .B1(_0943_));
 sg13g2_o21ai_1 _3831_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0944_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[36] ),
    .A2(net643));
 sg13g2_a21oi_1 _3832_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2210_),
    .A2(net642),
    .Y(_0135_),
    .B1(_0944_));
 sg13g2_o21ai_1 _3833_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0945_),
    .VSS(VGND),
    .A1(net481),
    .A2(net664));
 sg13g2_a21oi_1 _3834_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2209_),
    .A2(net664),
    .Y(_0136_),
    .B1(_0945_));
 sg13g2_o21ai_1 _3835_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0946_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[38] ),
    .A2(net643));
 sg13g2_a21oi_1 _3836_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2209_),
    .A2(net643),
    .Y(_0137_),
    .B1(_0946_));
 sg13g2_o21ai_1 _3837_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0947_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[38] ),
    .A2(net656));
 sg13g2_a21oi_1 _3838_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2208_),
    .A2(net656),
    .Y(_0138_),
    .B1(_0947_));
 sg13g2_o21ai_1 _3839_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0948_),
    .VSS(VGND),
    .A1(net422),
    .A2(net656));
 sg13g2_a21oi_1 _3840_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2207_),
    .A2(net653),
    .Y(_0139_),
    .B1(_0948_));
 sg13g2_o21ai_1 _3841_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0949_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .A2(net642));
 sg13g2_a21oi_1 _3842_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2207_),
    .A2(net641),
    .Y(_0140_),
    .B1(_0949_));
 sg13g2_o21ai_1 _3843_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0950_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .A2(net656));
 sg13g2_a21oi_1 _3844_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2206_),
    .A2(net656),
    .Y(_0141_),
    .B1(_0950_));
 sg13g2_o21ai_1 _3845_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0951_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[42] ),
    .A2(net665));
 sg13g2_a21oi_1 _3846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2205_),
    .A2(net665),
    .Y(_0142_),
    .B1(_0951_));
 sg13g2_o21ai_1 _3847_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0952_),
    .VSS(VGND),
    .A1(net860),
    .A2(net643));
 sg13g2_a21oi_1 _3848_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2205_),
    .A2(net643),
    .Y(_0143_),
    .B1(_0952_));
 sg13g2_o21ai_1 _3849_ (.B1(net831),
    .VDD(VPWR),
    .Y(_0953_),
    .VSS(VGND),
    .A1(net860),
    .A2(net664));
 sg13g2_a21oi_1 _3850_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2204_),
    .A2(net664),
    .Y(_0144_),
    .B1(_0953_));
 sg13g2_o21ai_1 _3851_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0954_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[45] ),
    .A2(net657));
 sg13g2_a21oi_1 _3852_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2203_),
    .A2(net657),
    .Y(_0145_),
    .B1(_0954_));
 sg13g2_o21ai_1 _3853_ (.B1(net826),
    .VDD(VPWR),
    .Y(_0955_),
    .VSS(VGND),
    .A1(net530),
    .A2(net658));
 sg13g2_a21oi_1 _3854_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2202_),
    .A2(net658),
    .Y(_0146_),
    .B1(_0955_));
 sg13g2_o21ai_1 _3855_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0956_),
    .VSS(VGND),
    .A1(net1008),
    .A2(net642));
 sg13g2_a21oi_1 _3856_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2202_),
    .A2(net642),
    .Y(_0147_),
    .B1(_0956_));
 sg13g2_o21ai_1 _3857_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0957_),
    .VSS(VGND),
    .A1(net1008),
    .A2(net658));
 sg13g2_a21oi_1 _3858_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2201_),
    .A2(net658),
    .Y(_0148_),
    .B1(_0957_));
 sg13g2_o21ai_1 _3859_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0958_),
    .VSS(VGND),
    .A1(net434),
    .A2(net664));
 sg13g2_a21oi_1 _3860_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2200_),
    .A2(net664),
    .Y(_0149_),
    .B1(_0958_));
 sg13g2_o21ai_1 _3861_ (.B1(net831),
    .VDD(VPWR),
    .Y(_0959_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .A2(net643));
 sg13g2_a21oi_1 _3862_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2200_),
    .A2(net645),
    .Y(_0150_),
    .B1(_0959_));
 sg13g2_o21ai_1 _3863_ (.B1(net830),
    .VDD(VPWR),
    .Y(_0960_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .A2(net665));
 sg13g2_a21oi_1 _3864_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2199_),
    .A2(net665),
    .Y(_0151_),
    .B1(_0960_));
 sg13g2_o21ai_1 _3865_ (.B1(net829),
    .VDD(VPWR),
    .Y(_0961_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[52] ),
    .A2(net665));
 sg13g2_a21oi_1 _3866_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2198_),
    .A2(net657),
    .Y(_0152_),
    .B1(_0961_));
 sg13g2_o21ai_1 _3867_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0962_),
    .VSS(VGND),
    .A1(net443),
    .A2(net657));
 sg13g2_a21oi_1 _3868_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2197_),
    .A2(net657),
    .Y(_0153_),
    .B1(_0962_));
 sg13g2_o21ai_1 _3869_ (.B1(net825),
    .VDD(VPWR),
    .Y(_0963_),
    .VSS(VGND),
    .A1(net398),
    .A2(net645));
 sg13g2_a21oi_1 _3870_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2197_),
    .A2(net645),
    .Y(_0154_),
    .B1(_0963_));
 sg13g2_o21ai_1 _3871_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0964_),
    .VSS(VGND),
    .A1(net398),
    .A2(net665));
 sg13g2_a21oi_1 _3872_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2196_),
    .A2(net671),
    .Y(_0155_),
    .B1(_0964_));
 sg13g2_o21ai_1 _3873_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0965_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[57] ),
    .A2(net646));
 sg13g2_a21oi_1 _3874_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2196_),
    .A2(net646),
    .Y(_0156_),
    .B1(_0965_));
 sg13g2_o21ai_1 _3875_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0966_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[57] ),
    .A2(net671));
 sg13g2_a21oi_1 _3876_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2195_),
    .A2(net671),
    .Y(_0157_),
    .B1(_0966_));
 sg13g2_o21ai_1 _3877_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0967_),
    .VSS(VGND),
    .A1(net557),
    .A2(net670));
 sg13g2_a21oi_1 _3878_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2194_),
    .A2(net670),
    .Y(_0158_),
    .B1(_0967_));
 sg13g2_o21ai_1 _3879_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0968_),
    .VSS(VGND),
    .A1(net866),
    .A2(net676));
 sg13g2_a21oi_1 _3880_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2193_),
    .A2(net676),
    .Y(_0159_),
    .B1(_0968_));
 sg13g2_o21ai_1 _3881_ (.B1(net840),
    .VDD(VPWR),
    .Y(_0969_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[60] ),
    .A2(net677));
 sg13g2_a21oi_1 _3882_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2192_),
    .A2(net676),
    .Y(_0160_),
    .B1(_0969_));
 sg13g2_o21ai_1 _3883_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0970_),
    .VSS(VGND),
    .A1(net474),
    .A2(net649));
 sg13g2_a21oi_1 _3884_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2192_),
    .A2(net649),
    .Y(_0161_),
    .B1(_0970_));
 sg13g2_o21ai_1 _3885_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0971_),
    .VSS(VGND),
    .A1(net474),
    .A2(net670));
 sg13g2_a21oi_1 _3886_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2191_),
    .A2(net670),
    .Y(_0162_),
    .B1(_0971_));
 sg13g2_o21ai_1 _3887_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0972_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[63] ),
    .A2(net671));
 sg13g2_a21oi_1 _3888_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2190_),
    .A2(net671),
    .Y(_0163_),
    .B1(_0972_));
 sg13g2_o21ai_1 _3889_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0973_),
    .VSS(VGND),
    .A1(net522),
    .A2(net647));
 sg13g2_a21oi_1 _3890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2190_),
    .A2(net647),
    .Y(_0164_),
    .B1(_0973_));
 sg13g2_o21ai_1 _3891_ (.B1(net835),
    .VDD(VPWR),
    .Y(_0974_),
    .VSS(VGND),
    .A1(net522),
    .A2(net669));
 sg13g2_a21oi_1 _3892_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2189_),
    .A2(net669),
    .Y(_0165_),
    .B1(_0974_));
 sg13g2_o21ai_1 _3893_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0975_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[66] ),
    .A2(net676));
 sg13g2_a21oi_1 _3894_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2188_),
    .A2(net676),
    .Y(_0166_),
    .B1(_0975_));
 sg13g2_o21ai_1 _3895_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0976_),
    .VSS(VGND),
    .A1(net889),
    .A2(net676));
 sg13g2_a21oi_1 _3896_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2187_),
    .A2(net678),
    .Y(_0167_),
    .B1(_0976_));
 sg13g2_o21ai_1 _3897_ (.B1(net840),
    .VDD(VPWR),
    .Y(_0977_),
    .VSS(VGND),
    .A1(net962),
    .A2(net649));
 sg13g2_a21oi_1 _3898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2187_),
    .A2(net649),
    .Y(_0168_),
    .B1(_0977_));
 sg13g2_o21ai_1 _3899_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0978_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .A2(net676));
 sg13g2_a21oi_1 _3900_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2186_),
    .A2(net670),
    .Y(_0169_),
    .B1(_0978_));
 sg13g2_o21ai_1 _3901_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0979_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[70] ),
    .A2(net669));
 sg13g2_a21oi_1 _3902_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2185_),
    .A2(net671),
    .Y(_0170_),
    .B1(_0979_));
 sg13g2_o21ai_1 _3903_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0980_),
    .VSS(VGND),
    .A1(net482),
    .A2(net646));
 sg13g2_a21oi_1 _3904_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2185_),
    .A2(net647),
    .Y(_0171_),
    .B1(_0980_));
 sg13g2_o21ai_1 _3905_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0981_),
    .VSS(VGND),
    .A1(net482),
    .A2(net669));
 sg13g2_a21oi_1 _3906_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2184_),
    .A2(net670),
    .Y(_0172_),
    .B1(_0981_));
 sg13g2_o21ai_1 _3907_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0982_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[73] ),
    .A2(net678));
 sg13g2_a21oi_1 _3908_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2183_),
    .A2(net678),
    .Y(_0173_),
    .B1(_0982_));
 sg13g2_o21ai_1 _3909_ (.B1(net840),
    .VDD(VPWR),
    .Y(_0983_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[74] ),
    .A2(net678));
 sg13g2_a21oi_1 _3910_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2182_),
    .A2(net678),
    .Y(_0174_),
    .B1(_0983_));
 sg13g2_o21ai_1 _3911_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0984_),
    .VSS(VGND),
    .A1(net404),
    .A2(net649));
 sg13g2_a21oi_1 _3912_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2182_),
    .A2(net649),
    .Y(_0175_),
    .B1(_0984_));
 sg13g2_o21ai_1 _3913_ (.B1(net839),
    .VDD(VPWR),
    .Y(_0985_),
    .VSS(VGND),
    .A1(net404),
    .A2(net676));
 sg13g2_a21oi_1 _3914_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2181_),
    .A2(net670),
    .Y(_0176_),
    .B1(_0985_));
 sg13g2_o21ai_1 _3915_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0986_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[77] ),
    .A2(net669));
 sg13g2_a21oi_1 _3916_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2180_),
    .A2(net669),
    .Y(_0177_),
    .B1(_0986_));
 sg13g2_o21ai_1 _3917_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0987_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[78] ),
    .A2(net669));
 sg13g2_a21oi_1 _3918_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2179_),
    .A2(net669),
    .Y(_0178_),
    .B1(_0987_));
 sg13g2_o21ai_1 _3919_ (.B1(net834),
    .VDD(VPWR),
    .Y(_0988_),
    .VSS(VGND),
    .A1(net886),
    .A2(net647));
 sg13g2_a21oi_1 _3920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2179_),
    .A2(net647),
    .Y(_0179_),
    .B1(_0988_));
 sg13g2_o21ai_1 _3921_ (.B1(net840),
    .VDD(VPWR),
    .Y(_0989_),
    .VSS(VGND),
    .A1(net886),
    .A2(net677));
 sg13g2_a21oi_1 _3922_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2177_),
    .A2(net677),
    .Y(_0180_),
    .B1(_0989_));
 sg13g2_o21ai_1 _3923_ (.B1(net840),
    .VDD(VPWR),
    .Y(_0990_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[81] ),
    .A2(net677));
 sg13g2_a21oi_1 _3924_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2176_),
    .A2(net677),
    .Y(_0181_),
    .B1(_0990_));
 sg13g2_o21ai_1 _3925_ (.B1(net841),
    .VDD(VPWR),
    .Y(_0991_),
    .VSS(VGND),
    .A1(net930),
    .A2(net649));
 sg13g2_a21oi_1 _3926_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2176_),
    .A2(net650),
    .Y(_0182_),
    .B1(_0991_));
 sg13g2_o21ai_1 _3927_ (.B1(net841),
    .VDD(VPWR),
    .Y(_0992_),
    .VSS(VGND),
    .A1(net930),
    .A2(net674));
 sg13g2_a21oi_1 _3928_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2175_),
    .A2(net674),
    .Y(_0183_),
    .B1(_0992_));
 sg13g2_o21ai_1 _3929_ (.B1(net837),
    .VDD(VPWR),
    .Y(_0993_),
    .VSS(VGND),
    .A1(net878),
    .A2(net673));
 sg13g2_a21oi_1 _3930_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2174_),
    .A2(net673),
    .Y(_0184_),
    .B1(_0993_));
 sg13g2_o21ai_1 _3931_ (.B1(net837),
    .VDD(VPWR),
    .Y(_0994_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .A2(net650));
 sg13g2_a21oi_1 _3932_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2174_),
    .A2(net650),
    .Y(_0185_),
    .B1(_0994_));
 sg13g2_o21ai_1 _3933_ (.B1(net838),
    .VDD(VPWR),
    .Y(_0995_),
    .VSS(VGND),
    .A1(net544),
    .A2(net675));
 sg13g2_a21oi_1 _3934_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2173_),
    .A2(net675),
    .Y(_0186_),
    .B1(_0995_));
 sg13g2_o21ai_1 _3935_ (.B1(net836),
    .VDD(VPWR),
    .Y(_0996_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .A2(net646));
 sg13g2_a21oi_1 _3936_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2173_),
    .A2(net646),
    .Y(_0187_),
    .B1(_0996_));
 sg13g2_o21ai_1 _3937_ (.B1(net836),
    .VDD(VPWR),
    .Y(_0997_),
    .VSS(VGND),
    .A1(net541),
    .A2(net668));
 sg13g2_a21oi_1 _3938_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2172_),
    .A2(net667),
    .Y(_0188_),
    .B1(_0997_));
 sg13g2_o21ai_1 _3939_ (.B1(net836),
    .VDD(VPWR),
    .Y(_0998_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .A2(net646));
 sg13g2_a21oi_1 _3940_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2172_),
    .A2(net646),
    .Y(_0189_),
    .B1(_0998_));
 sg13g2_o21ai_1 _3941_ (.B1(net838),
    .VDD(VPWR),
    .Y(_0999_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .A2(net672));
 sg13g2_a21oi_1 _3942_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2171_),
    .A2(net672),
    .Y(_0190_),
    .B1(_0999_));
 sg13g2_o21ai_1 _3943_ (.B1(net837),
    .VDD(VPWR),
    .Y(_1000_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[91] ),
    .A2(net673));
 sg13g2_a21oi_1 _3944_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2170_),
    .A2(net673),
    .Y(_0191_),
    .B1(_1000_));
 sg13g2_o21ai_1 _3945_ (.B1(net837),
    .VDD(VPWR),
    .Y(_1001_),
    .VSS(VGND),
    .A1(net401),
    .A2(net648));
 sg13g2_a21oi_1 _3946_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2170_),
    .A2(net648),
    .Y(_0192_),
    .B1(_1001_));
 sg13g2_o21ai_1 _3947_ (.B1(net838),
    .VDD(VPWR),
    .Y(_1002_),
    .VSS(VGND),
    .A1(net401),
    .A2(net672));
 sg13g2_a21oi_1 _3948_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2169_),
    .A2(net672),
    .Y(_0193_),
    .B1(_1002_));
 sg13g2_o21ai_1 _3949_ (.B1(net840),
    .VDD(VPWR),
    .Y(_1003_),
    .VSS(VGND),
    .A1(net867),
    .A2(net674));
 sg13g2_a21oi_1 _3950_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2168_),
    .A2(net677),
    .Y(_0194_),
    .B1(_1003_));
 sg13g2_o21ai_1 _3951_ (.B1(net840),
    .VDD(VPWR),
    .Y(_1004_),
    .VSS(VGND),
    .A1(net556),
    .A2(net677));
 sg13g2_a21oi_1 _3952_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2167_),
    .A2(net677),
    .Y(_0195_),
    .B1(_1004_));
 sg13g2_o21ai_1 _3953_ (.B1(net841),
    .VDD(VPWR),
    .Y(_1005_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .A2(net648));
 sg13g2_a21oi_1 _3954_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2167_),
    .A2(net649),
    .Y(_0196_),
    .B1(_1005_));
 sg13g2_o21ai_1 _3955_ (.B1(net841),
    .VDD(VPWR),
    .Y(_1006_),
    .VSS(VGND),
    .A1(net961),
    .A2(net674));
 sg13g2_a21oi_1 _3956_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2166_),
    .A2(net674),
    .Y(_0197_),
    .B1(_1006_));
 sg13g2_o21ai_1 _3957_ (.B1(net837),
    .VDD(VPWR),
    .Y(_1007_),
    .VSS(VGND),
    .A1(net562),
    .A2(net674));
 sg13g2_a21oi_1 _3958_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2165_),
    .A2(net674),
    .Y(_0198_),
    .B1(_1007_));
 sg13g2_o21ai_1 _3959_ (.B1(net837),
    .VDD(VPWR),
    .Y(_1008_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .A2(net648));
 sg13g2_a21oi_1 _3960_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2165_),
    .A2(net650),
    .Y(_0199_),
    .B1(_1008_));
 sg13g2_o21ai_1 _3961_ (.B1(net838),
    .VDD(VPWR),
    .Y(_1009_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .A2(net672));
 sg13g2_a21oi_1 _3962_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2164_),
    .A2(net672),
    .Y(_0200_),
    .B1(_1009_));
 sg13g2_o21ai_1 _3963_ (.B1(net836),
    .VDD(VPWR),
    .Y(_1010_),
    .VSS(VGND),
    .A1(net500),
    .A2(net667));
 sg13g2_a21oi_1 _3964_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2163_),
    .A2(net668),
    .Y(_0201_),
    .B1(_1010_));
 sg13g2_o21ai_1 _3965_ (.B1(net836),
    .VDD(VPWR),
    .Y(_1011_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[102] ),
    .A2(net667));
 sg13g2_a21oi_1 _3966_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2162_),
    .A2(net667),
    .Y(_0202_),
    .B1(_1011_));
 sg13g2_o21ai_1 _3967_ (.B1(net838),
    .VDD(VPWR),
    .Y(_1012_),
    .VSS(VGND),
    .A1(net454),
    .A2(net648));
 sg13g2_a21oi_1 _3968_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2162_),
    .A2(net648),
    .Y(_0203_),
    .B1(_1012_));
 sg13g2_o21ai_1 _3969_ (.B1(net841),
    .VDD(VPWR),
    .Y(_1013_),
    .VSS(VGND),
    .A1(net454),
    .A2(net673));
 sg13g2_a21oi_1 _3970_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2161_),
    .A2(net673),
    .Y(_0204_),
    .B1(_1013_));
 sg13g2_o21ai_1 _3971_ (.B1(net837),
    .VDD(VPWR),
    .Y(_1014_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[105] ),
    .A2(net673));
 sg13g2_a21oi_1 _3972_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2160_),
    .A2(net673),
    .Y(_0205_),
    .B1(_1014_));
 sg13g2_o21ai_1 _3973_ (.B1(net837),
    .VDD(VPWR),
    .Y(_1015_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[106] ),
    .A2(net672));
 sg13g2_a21oi_1 _3974_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2159_),
    .A2(net672),
    .Y(_0206_),
    .B1(_1015_));
 sg13g2_o21ai_1 _3975_ (.B1(net838),
    .VDD(VPWR),
    .Y(_1016_),
    .VSS(VGND),
    .A1(net540),
    .A2(net648));
 sg13g2_a21oi_1 _3976_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2159_),
    .A2(net648),
    .Y(_0207_),
    .B1(_1016_));
 sg13g2_o21ai_1 _3977_ (.B1(net838),
    .VDD(VPWR),
    .Y(_1017_),
    .VSS(VGND),
    .A1(\ppwm_i.u_ppwm.u_mem.memory[108] ),
    .A2(net667));
 sg13g2_a21oi_1 _3978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2158_),
    .A2(net667),
    .Y(_0208_),
    .B1(_1017_));
 sg13g2_o21ai_1 _3979_ (.B1(net836),
    .VDD(VPWR),
    .Y(_1018_),
    .VSS(VGND),
    .A1(net461),
    .A2(net667));
 sg13g2_a21oi_1 _3980_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2157_),
    .A2(net667),
    .Y(_0209_),
    .B1(_1018_));
 sg13g2_o21ai_1 _3981_ (.B1(net836),
    .VDD(VPWR),
    .Y(_1019_),
    .VSS(VGND),
    .A1(net559),
    .A2(net668));
 sg13g2_a21oi_1 _3982_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2156_),
    .A2(net668),
    .Y(_0210_),
    .B1(_1019_));
 sg13g2_o21ai_1 _3983_ (.B1(net808),
    .VDD(VPWR),
    .Y(_1020_),
    .VSS(VGND),
    .A1(net971),
    .A2(net652));
 sg13g2_a21oi_1 _3984_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2156_),
    .A2(net646),
    .Y(_0211_),
    .B1(_1020_));
 sg13g2_nand2_2 _3985_ (.Y(_1021_),
    .A(net934),
    .B(_0906_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _3986_ (.Y(_1022_),
    .A(net652),
    .B(_1021_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3987_ (.B1(net808),
    .VDD(VPWR),
    .Y(_1023_),
    .VSS(VGND),
    .A1(net378),
    .A2(net680));
 sg13g2_a21oi_1 _3988_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net378),
    .A2(_1022_),
    .Y(_0212_),
    .B1(_1023_));
 sg13g2_nand3_1 _3989_ (.B(net652),
    .C(_1021_),
    .A(net1152),
    .Y(_1024_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _3990_ (.A(net1152),
    .B(net378),
    .X(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3991_ (.B1(net680),
    .VDD(VPWR),
    .Y(_1026_),
    .VSS(VGND),
    .A1(net1152),
    .A2(net378));
 sg13g2_o21ai_1 _3992_ (.B1(_1024_),
    .VDD(VPWR),
    .Y(_1027_),
    .VSS(VGND),
    .A1(_1025_),
    .A2(_1026_));
 sg13g2_and2_1 _3993_ (.A(net808),
    .B(_1027_),
    .X(_0213_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _3994_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net1051),
    .A2(_1021_),
    .Y(_1028_),
    .B1(net680));
 sg13g2_nand2_1 _3995_ (.Y(_1029_),
    .A(net1051),
    .B(_1025_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _3996_ (.A(net652),
    .B(_1029_),
    .Y(_1030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3997_ (.B1(net808),
    .VDD(VPWR),
    .Y(_1031_),
    .VSS(VGND),
    .A1(net1051),
    .A2(_1025_));
 sg13g2_nor3_1 _3998_ (.A(net1052),
    .B(_1030_),
    .C(_1031_),
    .Y(_0214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _3999_ (.B1(net1186),
    .VDD(VPWR),
    .Y(_1032_),
    .VSS(VGND),
    .A1(net883),
    .A2(_1021_));
 sg13g2_nand2b_1 _4000_ (.Y(_1033_),
    .B(_1032_),
    .A_N(_1030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4001_ (.Y(_1034_),
    .A(net1186),
    .B(_1030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4002_ (.X(_0215_),
    .A(net808),
    .B(_1033_),
    .C(_1034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4003_ (.B1(net1010),
    .VDD(VPWR),
    .Y(_1035_),
    .VSS(VGND),
    .A1(net883),
    .A2(_1021_));
 sg13g2_nand3_1 _4004_ (.B(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .C(_1030_),
    .A(net1010),
    .Y(_1036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4005_ (.Y(_1037_),
    .A(net807),
    .B(_1036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4006_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1034_),
    .A2(net1011),
    .Y(_0216_),
    .B1(_1037_));
 sg13g2_nand3_1 _4007_ (.B(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .C(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .A(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .Y(_1038_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4008_ (.B1(net883),
    .VDD(VPWR),
    .Y(_1039_),
    .VSS(VGND),
    .A1(_1029_),
    .A2(_1038_));
 sg13g2_a21oi_1 _4009_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1022_),
    .A2(_1039_),
    .Y(_1040_),
    .B1(net796));
 sg13g2_nand2b_1 _4010_ (.Y(_1041_),
    .B(_1036_),
    .A_N(net1155),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4011_ (.A(_1040_),
    .B(net1156),
    .X(_0217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4012_ (.Y(_1042_),
    .A(net512),
    .B(_1040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _4013_ (.B(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .C(net806),
    .Y(_1043_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net512));
 sg13g2_o21ai_1 _4014_ (.B1(net513),
    .VDD(VPWR),
    .Y(_0218_),
    .VSS(VGND),
    .A1(_1036_),
    .A2(_1043_));
 sg13g2_nor3_1 _4015_ (.A(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .B(_0397_),
    .C(_1034_),
    .Y(_1044_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4016_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net934),
    .A2(_0906_),
    .Y(_1045_),
    .B1(net883));
 sg13g2_nor3_1 _4017_ (.A(net796),
    .B(_1044_),
    .C(net935),
    .Y(_0219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4018_ (.A(net2),
    .B_N(net1),
    .Y(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4019_ (.B1(net805),
    .VDD(VPWR),
    .Y(_1047_),
    .VSS(VGND),
    .A1(\falu_i.falutop.i2c_inst.state[0] ),
    .A2(_1046_));
 sg13g2_nor2_1 _4020_ (.A(net459),
    .B(_1047_),
    .Y(_0220_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _4021_ (.A(\falu_i.falutop.i2c_inst.state[0] ),
    .B_N(net459),
    .Y(_1048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4022_ (.A(_2433_),
    .B(_1048_),
    .Y(_1049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4023_ (.A(net1),
    .B(_1049_),
    .X(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4024_ (.Y(_1051_),
    .A(net2),
    .B(_1050_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4025_ (.Y(_1052_),
    .A(net1013),
    .B(_2438_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4026_ (.B1(_1051_),
    .VDD(VPWR),
    .Y(_1053_),
    .VSS(VGND),
    .A1(_1049_),
    .A2(_1052_));
 sg13g2_mux2_1 _4027_ (.A0(net459),
    .A1(net1015),
    .S(_2442_),
    .X(_1054_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4028_ (.B1(net816),
    .VDD(VPWR),
    .Y(_1055_),
    .VSS(VGND),
    .A1(net459),
    .A2(_1053_));
 sg13g2_nor2_1 _4029_ (.A(_1054_),
    .B(_1055_),
    .Y(_0221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4030_ (.A(net1043),
    .B(_1049_),
    .Y(_1056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4031_ (.A(net459),
    .B(net1015),
    .Y(_1057_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4032_ (.Y(_1058_),
    .A(_2442_),
    .B(_0901_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4033_ (.Y(_1059_),
    .B(_1058_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1057_));
 sg13g2_nor2_1 _4034_ (.A(_1050_),
    .B(_1056_),
    .Y(_1060_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4035_ (.B1(net804),
    .VDD(VPWR),
    .Y(_1061_),
    .VSS(VGND),
    .A1(net1043),
    .A2(_1059_));
 sg13g2_a21oi_1 _4036_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1059_),
    .A2(_1060_),
    .Y(_0222_),
    .B1(_1061_));
 sg13g2_nor3_1 _4037_ (.A(_2445_),
    .B(_0343_),
    .C(_1049_),
    .Y(_1062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4038_ (.A(_1050_),
    .B(_1062_),
    .Y(_1063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4039_ (.B1(net816),
    .VDD(VPWR),
    .Y(_1064_),
    .VSS(VGND),
    .A1(net1028),
    .A2(_1059_));
 sg13g2_a21oi_1 _4040_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1059_),
    .A2(_1063_),
    .Y(_0223_),
    .B1(_1064_));
 sg13g2_nand2b_1 _4041_ (.Y(_1065_),
    .B(_1059_),
    .A_N(_1053_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4042_ (.B1(_1065_),
    .VDD(VPWR),
    .Y(_1066_),
    .VSS(VGND),
    .A1(net1006),
    .A2(_1059_));
 sg13g2_nor2_1 _4043_ (.A(net797),
    .B(_1066_),
    .Y(_0224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4044_ (.Y(_1067_),
    .B(_2441_),
    .A_N(_1049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4045_ (.Y(_1068_),
    .A(_1051_),
    .B(_1067_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4046_ (.B1(_1059_),
    .VDD(VPWR),
    .Y(_1069_),
    .VSS(VGND),
    .A1(_2440_),
    .A2(_1057_));
 sg13g2_a22oi_1 _4047_ (.Y(_1070_),
    .B1(_1069_),
    .B2(net985),
    .A2(_1068_),
    .A1(_1059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4048_ (.A(net797),
    .B(_1070_),
    .Y(_0225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4049_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2441_),
    .A2(_0901_),
    .Y(_1071_),
    .B1(_1057_));
 sg13g2_a22oi_1 _4050_ (.Y(_1072_),
    .B1(_1071_),
    .B2(net1016),
    .A2(_1057_),
    .A1(_1046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4051_ (.A(net797),
    .B(_1072_),
    .Y(_0226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _4052_ (.A(_2291_),
    .B(\falu_i.falutop.i2c_inst.op[1] ),
    .C(_2292_),
    .D(_2293_),
    .Y(_1073_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or4_1 _4053_ (.A(_2291_),
    .B(\falu_i.falutop.i2c_inst.op[1] ),
    .C(_2292_),
    .D(_2293_),
    .X(_1074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4054_ (.A(net380),
    .B(_1074_),
    .Y(_1075_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4055_ (.Y(_1076_),
    .B(net639),
    .A_N(\falu_i.falutop.div_inst.done ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4056_ (.A(_2294_),
    .B(_1074_),
    .Y(_1077_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4057_ (.Y(_1078_),
    .A(net815),
    .B(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4058_ (.A(net380),
    .B(net622),
    .Y(_0227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4059_ (.A0(net848),
    .A1(\falu_i.falutop.data_in[0] ),
    .S(net684),
    .X(_0228_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4060_ (.A0(net901),
    .A1(\falu_i.falutop.data_in[1] ),
    .S(net684),
    .X(_0229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4061_ (.A0(net972),
    .A1(\falu_i.falutop.data_in[2] ),
    .S(net685),
    .X(_0230_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4062_ (.A0(net992),
    .A1(\falu_i.falutop.data_in[3] ),
    .S(net685),
    .X(_0231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4063_ (.A0(net881),
    .A1(\falu_i.falutop.data_in[4] ),
    .S(net685),
    .X(_0232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4064_ (.A0(net869),
    .A1(\falu_i.falutop.data_in[5] ),
    .S(net684),
    .X(_0233_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4065_ (.A0(net850),
    .A1(\falu_i.falutop.data_in[6] ),
    .S(net684),
    .X(_0234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4066_ (.A0(net871),
    .A1(net777),
    .S(net684),
    .X(_0235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4067_ (.A0(net873),
    .A1(\falu_i.falutop.data_in[8] ),
    .S(net684),
    .X(_0236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4068_ (.A0(net899),
    .A1(\falu_i.falutop.data_in[9] ),
    .S(net685),
    .X(_0237_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4069_ (.A0(net945),
    .A1(\falu_i.falutop.data_in[10] ),
    .S(net685),
    .X(_0238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4070_ (.A0(net858),
    .A1(\falu_i.falutop.data_in[11] ),
    .S(net685),
    .X(_0239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4071_ (.A0(net926),
    .A1(\falu_i.falutop.data_in[12] ),
    .S(net685),
    .X(_0240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4072_ (.A0(net894),
    .A1(\falu_i.falutop.data_in[13] ),
    .S(net684),
    .X(_0241_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4073_ (.A0(net861),
    .A1(\falu_i.falutop.data_in[14] ),
    .S(net687),
    .X(_0242_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4074_ (.A0(net908),
    .A1(net775),
    .S(net684),
    .X(_0243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4075_ (.A(\falu_i.falutop.i2c_inst.result[10] ),
    .B(_0343_),
    .X(_1079_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4076_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(\falu_i.falutop.i2c_inst.result[9] ),
    .A2(_2445_),
    .Y(_1080_),
    .B1(\falu_i.falutop.i2c_inst.counter[2] ));
 sg13g2_a221oi_1 _4077_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\falu_i.falutop.i2c_inst.result[8] ),
    .C1(_1079_),
    .B1(_2438_),
    .A1(\falu_i.falutop.i2c_inst.result[11] ),
    .Y(_1081_),
    .A2(_2432_));
 sg13g2_a22oi_1 _4078_ (.Y(_1082_),
    .B1(_2438_),
    .B2(\falu_i.falutop.i2c_inst.result[12] ),
    .A2(_2432_),
    .A1(\falu_i.falutop.i2c_inst.result[15] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4079_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(\falu_i.falutop.i2c_inst.result[14] ),
    .C1(_2154_),
    .B1(_0343_),
    .A1(\falu_i.falutop.i2c_inst.result[13] ),
    .Y(_1083_),
    .A2(_2445_));
 sg13g2_a22oi_1 _4080_ (.Y(_1084_),
    .B1(_1082_),
    .B2(_1083_),
    .A2(_1081_),
    .A1(_1080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4081_ (.Y(_1085_),
    .B1(_2438_),
    .B2(\falu_i.falutop.i2c_inst.result[0] ),
    .A2(_2432_),
    .A1(\falu_i.falutop.i2c_inst.result[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4082_ (.Y(_1086_),
    .B1(_0343_),
    .B2(\falu_i.falutop.i2c_inst.result[2] ),
    .A2(_2445_),
    .A1(\falu_i.falutop.i2c_inst.result[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4083_ (.Y(_1087_),
    .A(_1085_),
    .B(_1086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4084_ (.Y(_1088_),
    .A(_2430_),
    .B(_1087_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4085_ (.Y(_1089_),
    .B1(_2438_),
    .B2(\falu_i.falutop.i2c_inst.result[4] ),
    .A2(_2432_),
    .A1(\falu_i.falutop.i2c_inst.result[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4086_ (.Y(_1090_),
    .B1(_0343_),
    .B2(\falu_i.falutop.i2c_inst.result[6] ),
    .A2(_2445_),
    .A1(\falu_i.falutop.i2c_inst.result[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4087_ (.Y(_1091_),
    .A(_1089_),
    .B(_1090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4088_ (.Y(_1092_),
    .A(_1048_),
    .B(_1088_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4089_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net986),
    .C1(_1092_),
    .B1(_1091_),
    .A1(net985),
    .Y(_1093_),
    .A2(_1084_));
 sg13g2_o21ai_1 _4090_ (.B1(net805),
    .VDD(VPWR),
    .Y(_1094_),
    .VSS(VGND),
    .A1(net996),
    .A2(_1048_));
 sg13g2_nor2_1 _4091_ (.A(_1093_),
    .B(net997),
    .Y(_0244_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4092_ (.B(\falu_i.falutop.div_inst.i[1] ),
    .C(net525),
    .A(net409),
    .Y(_1095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4093_ (.Y(_1096_),
    .B(\falu_i.falutop.div_inst.busy ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net778));
 sg13g2_nor2b_2 _4094_ (.A(_1096_),
    .B_N(_1095_),
    .Y(_1097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4095_ (.Y(_1098_),
    .B(_1095_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1096_));
 sg13g2_nor4_1 _4096_ (.A(net983),
    .B(net999),
    .C(net1054),
    .D(net920),
    .Y(_1099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _4097_ (.A(net413),
    .B(net1081),
    .C(net967),
    .D(net891),
    .Y(_1100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4098_ (.Y(_1101_),
    .A(_1099_),
    .B(_1100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4099_ (.VDD(VPWR),
    .Y(_1102_),
    .A(_1101_),
    .VSS(VGND));
 sg13g2_and2_1 _4100_ (.A(net778),
    .B(_1101_),
    .X(_1103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4101_ (.Y(_1104_),
    .A(net778),
    .B(_1101_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4102_ (.A(_1097_),
    .B(_1103_),
    .Y(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4103_ (.Y(_1106_),
    .A(_1098_),
    .B(_1104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4104_ (.A(net779),
    .B_N(net396),
    .Y(_1107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4105_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net779),
    .A2(net952),
    .Y(_1108_),
    .B1(_1107_));
 sg13g2_nor2_1 _4106_ (.A(net1009),
    .B(net606),
    .Y(_1109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4107_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net606),
    .A2(_1108_),
    .Y(_0245_),
    .B1(_1109_));
 sg13g2_xor2_1 _4108_ (.B(\falu_i.falutop.div_inst.acc[7] ),
    .A(\falu_i.falutop.div_inst.b1[7] ),
    .X(_1110_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4109_ (.A(\falu_i.falutop.div_inst.b1[6] ),
    .B_N(\falu_i.falutop.div_inst.acc[6] ),
    .Y(_1111_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4110_ (.A(\falu_i.falutop.div_inst.b1[5] ),
    .B_N(\falu_i.falutop.div_inst.acc[5] ),
    .Y(_1112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4111_ (.A(\falu_i.falutop.div_inst.b1[4] ),
    .B_N(\falu_i.falutop.div_inst.acc[4] ),
    .Y(_1113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4112_ (.A(\falu_i.falutop.div_inst.b1[3] ),
    .B_N(\falu_i.falutop.div_inst.acc[3] ),
    .Y(_1114_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4113_ (.A(\falu_i.falutop.div_inst.b1[2] ),
    .B_N(\falu_i.falutop.div_inst.acc[2] ),
    .Y(_1115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4114_ (.Y(_1116_),
    .B(\falu_i.falutop.div_inst.acc[1] ),
    .A_N(\falu_i.falutop.div_inst.b1[1] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4115_ (.A(\falu_i.falutop.div_inst.acc[0] ),
    .B_N(\falu_i.falutop.div_inst.b1[0] ),
    .Y(_1117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4116_ (.B(\falu_i.falutop.div_inst.acc[1] ),
    .A(\falu_i.falutop.div_inst.b1[1] ),
    .X(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4117_ (.B1(_1116_),
    .VDD(VPWR),
    .Y(_1119_),
    .VSS(VGND),
    .A1(_1117_),
    .A2(_1118_));
 sg13g2_xnor2_1 _4118_ (.Y(_1120_),
    .A(\falu_i.falutop.div_inst.b1[2] ),
    .B(\falu_i.falutop.div_inst.acc[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4119_ (.A2(_1120_),
    .A1(_1119_),
    .B1(_1115_),
    .X(_1121_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4120_ (.Y(_1122_),
    .A(\falu_i.falutop.div_inst.b1[3] ),
    .B(\falu_i.falutop.div_inst.acc[3] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4121_ (.A2(_1122_),
    .A1(_1121_),
    .B1(_1114_),
    .X(_1123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4122_ (.Y(_1124_),
    .A(\falu_i.falutop.div_inst.b1[4] ),
    .B(\falu_i.falutop.div_inst.acc[4] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4123_ (.A2(_1124_),
    .A1(_1123_),
    .B1(_1113_),
    .X(_1125_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4124_ (.Y(_1126_),
    .A(\falu_i.falutop.div_inst.b1[5] ),
    .B(\falu_i.falutop.div_inst.acc[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4125_ (.A2(_1126_),
    .A1(_1125_),
    .B1(_1112_),
    .X(_1127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4126_ (.Y(_1128_),
    .A(\falu_i.falutop.div_inst.b1[6] ),
    .B(\falu_i.falutop.div_inst.acc[6] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4127_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1127_),
    .A2(_1128_),
    .Y(_1129_),
    .B1(_1111_));
 sg13g2_nor2_1 _4128_ (.A(_1110_),
    .B(_1129_),
    .Y(_1130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4129_ (.A(net879),
    .B(_1130_),
    .Y(_1131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4130_ (.B1(_1131_),
    .VDD(VPWR),
    .Y(_1132_),
    .VSS(VGND),
    .A1(\falu_i.falutop.div_inst.b1[7] ),
    .A2(_2290_));
 sg13g2_a22oi_1 _4131_ (.Y(_1133_),
    .B1(net567),
    .B2(_1097_),
    .A2(net607),
    .A1(net910),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4132_ (.VDD(VPWR),
    .Y(_0246_),
    .A(net911),
    .VSS(VGND));
 sg13g2_nor2_2 _4133_ (.A(_1095_),
    .B(_1096_),
    .Y(_1134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4134_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net779),
    .A2(_1102_),
    .Y(_1135_),
    .B1(net633));
 sg13g2_nor2_1 _4135_ (.A(net797),
    .B(_1135_),
    .Y(_0247_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4136_ (.Y(_1136_),
    .A(net820),
    .B(_1074_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4137_ (.Y(_0248_),
    .B1(_2298_),
    .B2(net619),
    .A2(net833),
    .A1(_2291_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4138_ (.Y(_1137_),
    .B1(\falu_i.falutop.alu_inst.op[1] ),
    .B2(net619),
    .A2(net833),
    .A1(net1026),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4139_ (.VDD(VPWR),
    .Y(_0249_),
    .A(net1027),
    .VSS(VGND));
 sg13g2_a22oi_1 _4140_ (.Y(_0250_),
    .B1(_2299_),
    .B2(net619),
    .A2(net833),
    .A1(_2293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4141_ (.Y(_0251_),
    .B1(_2300_),
    .B2(net619),
    .A2(net833),
    .A1(_2292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4142_ (.A(net525),
    .B(\falu_i.falutop.div_inst.busy ),
    .X(_1138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4143_ (.Y(_1139_),
    .B(net525),
    .A_N(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4144_ (.Y(_0252_),
    .B1(net526),
    .B2(_1096_),
    .A2(_1138_),
    .A1(_1095_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4145_ (.Y(_1140_),
    .A(net917),
    .B(_1138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4146_ (.A(net409),
    .B(_1140_),
    .Y(_1141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4147_ (.A(net917),
    .B(_1138_),
    .Y(_1142_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4148_ (.A(net778),
    .B(_1141_),
    .C(net918),
    .Y(_0253_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4149_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2153_),
    .A2(_1140_),
    .Y(_0254_),
    .B1(net778));
 sg13g2_a22oi_1 _4150_ (.Y(_1143_),
    .B1(_1104_),
    .B2(net479),
    .A2(\falu_i.falutop.div_inst.b[0] ),
    .A1(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4151_ (.VDD(VPWR),
    .Y(_0255_),
    .A(net480),
    .VSS(VGND));
 sg13g2_mux2_1 _4152_ (.A0(net1005),
    .A1(net413),
    .S(_1103_),
    .X(_0256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4153_ (.A0(net1059),
    .A1(net891),
    .S(_1103_),
    .X(_0257_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4154_ (.Y(_1144_),
    .B1(_1104_),
    .B2(net994),
    .A2(net967),
    .A1(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4155_ (.VDD(VPWR),
    .Y(_0258_),
    .A(net995),
    .VSS(VGND));
 sg13g2_mux2_1 _4156_ (.A0(net1078),
    .A1(net999),
    .S(_1103_),
    .X(_0259_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4157_ (.A0(net1085),
    .A1(net983),
    .S(_1103_),
    .X(_0260_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4158_ (.A0(net1056),
    .A1(net920),
    .S(_1103_),
    .X(_0261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4159_ (.A0(\falu_i.falutop.div_inst.b1[7] ),
    .A1(net1054),
    .S(_1103_),
    .X(_0262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4160_ (.A(net797),
    .B(net607),
    .Y(_0263_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4161_ (.A(net568),
    .B_N(net633),
    .Y(_1145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4162_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1146_),
    .VSS(VGND),
    .A1(net1133),
    .A2(net634));
 sg13g2_nor2_1 _4163_ (.A(_1145_),
    .B(_1146_),
    .Y(_0264_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4164_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1147_),
    .VSS(VGND),
    .A1(net939),
    .A2(net635));
 sg13g2_a21oi_1 _4165_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2152_),
    .A2(net635),
    .Y(_0265_),
    .B1(net940));
 sg13g2_o21ai_1 _4166_ (.B1(net817),
    .VDD(VPWR),
    .Y(_1148_),
    .VSS(VGND),
    .A1(net978),
    .A2(net637));
 sg13g2_a21oi_1 _4167_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2151_),
    .A2(net637),
    .Y(_0266_),
    .B1(_1148_));
 sg13g2_o21ai_1 _4168_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1149_),
    .VSS(VGND),
    .A1(net947),
    .A2(net636));
 sg13g2_a21oi_1 _4169_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2150_),
    .A2(net636),
    .Y(_0267_),
    .B1(_1149_));
 sg13g2_o21ai_1 _4170_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1150_),
    .VSS(VGND),
    .A1(net905),
    .A2(net636));
 sg13g2_a21oi_1 _4171_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2149_),
    .A2(net636),
    .Y(_0268_),
    .B1(_1150_));
 sg13g2_o21ai_1 _4172_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1151_),
    .VSS(VGND),
    .A1(net937),
    .A2(net636));
 sg13g2_a21oi_1 _4173_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2148_),
    .A2(net636),
    .Y(_0269_),
    .B1(_1151_));
 sg13g2_o21ai_1 _4174_ (.B1(net819),
    .VDD(VPWR),
    .Y(_1152_),
    .VSS(VGND),
    .A1(net1037),
    .A2(net636));
 sg13g2_a21oi_1 _4175_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2147_),
    .A2(net637),
    .Y(_0270_),
    .B1(_1152_));
 sg13g2_o21ai_1 _4176_ (.B1(net819),
    .VDD(VPWR),
    .Y(_1153_),
    .VSS(VGND),
    .A1(\falu_i.falutop.div_inst.val[7] ),
    .A2(net637));
 sg13g2_a21oi_1 _4177_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2146_),
    .A2(net636),
    .Y(_0271_),
    .B1(_1153_));
 sg13g2_nand2_1 _4178_ (.Y(_1154_),
    .A(net479),
    .B(net568),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4179_ (.B(_1154_),
    .A(net1009),
    .X(_1155_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4180_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1156_),
    .VSS(VGND),
    .A1(net1116),
    .A2(net634));
 sg13g2_a21oi_1 _4181_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net634),
    .A2(_1155_),
    .Y(_0272_),
    .B1(_1156_));
 sg13g2_xnor2_1 _4182_ (.Y(_1157_),
    .A(_1117_),
    .B(_1118_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4183_ (.Y(_1158_),
    .A(net568),
    .B(_1157_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4184_ (.B1(_1158_),
    .VDD(VPWR),
    .Y(_1159_),
    .VSS(VGND),
    .A1(net498),
    .A2(net568));
 sg13g2_o21ai_1 _4185_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1160_),
    .VSS(VGND),
    .A1(net1098),
    .A2(net634));
 sg13g2_a21oi_1 _4186_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net634),
    .A2(_1159_),
    .Y(_0273_),
    .B1(_1160_));
 sg13g2_xnor2_1 _4187_ (.Y(_1161_),
    .A(_1119_),
    .B(_1120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4188_ (.Y(_1162_),
    .A(net568),
    .B(_1161_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4189_ (.B1(_1162_),
    .VDD(VPWR),
    .Y(_1163_),
    .VSS(VGND),
    .A1(net489),
    .A2(_1132_));
 sg13g2_o21ai_1 _4190_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1164_),
    .VSS(VGND),
    .A1(net1110),
    .A2(net634));
 sg13g2_a21oi_1 _4191_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1163_),
    .Y(_0274_),
    .B1(_1164_));
 sg13g2_xnor2_1 _4192_ (.Y(_1165_),
    .A(_1121_),
    .B(_1122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4193_ (.Y(_1166_),
    .A(net568),
    .B(_1165_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4194_ (.B1(_1166_),
    .VDD(VPWR),
    .Y(_1167_),
    .VSS(VGND),
    .A1(net494),
    .A2(net568));
 sg13g2_o21ai_1 _4195_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1168_),
    .VSS(VGND),
    .A1(net1119),
    .A2(net635));
 sg13g2_a21oi_1 _4196_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1167_),
    .Y(_0275_),
    .B1(_1168_));
 sg13g2_xnor2_1 _4197_ (.Y(_1169_),
    .A(_1123_),
    .B(_1124_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4198_ (.Y(_1170_),
    .A(net567),
    .B(_1169_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4199_ (.B1(_1170_),
    .VDD(VPWR),
    .Y(_1171_),
    .VSS(VGND),
    .A1(net856),
    .A2(net567));
 sg13g2_o21ai_1 _4200_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1172_),
    .VSS(VGND),
    .A1(net1124),
    .A2(net635));
 sg13g2_a21oi_1 _4201_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1171_),
    .Y(_0276_),
    .B1(_1172_));
 sg13g2_xnor2_1 _4202_ (.Y(_1173_),
    .A(_1125_),
    .B(_1126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4203_ (.Y(_1174_),
    .A(net567),
    .B(_1173_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4204_ (.B1(_1174_),
    .VDD(VPWR),
    .Y(_1175_),
    .VSS(VGND),
    .A1(net549),
    .A2(net567));
 sg13g2_o21ai_1 _4205_ (.B1(net803),
    .VDD(VPWR),
    .Y(_1176_),
    .VSS(VGND),
    .A1(net1106),
    .A2(net634));
 sg13g2_a21oi_1 _4206_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1175_),
    .Y(_0277_),
    .B1(_1176_));
 sg13g2_xnor2_1 _4207_ (.Y(_1177_),
    .A(_1127_),
    .B(_1128_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4208_ (.Y(_1178_),
    .A(net567),
    .B(_1177_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4209_ (.B1(_1178_),
    .VDD(VPWR),
    .Y(_1179_),
    .VSS(VGND),
    .A1(net931),
    .A2(net567));
 sg13g2_o21ai_1 _4210_ (.B1(net806),
    .VDD(VPWR),
    .Y(_1180_),
    .VSS(VGND),
    .A1(net1100),
    .A2(net633));
 sg13g2_a21oi_1 _4211_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net633),
    .A2(_1179_),
    .Y(_0278_),
    .B1(_1180_));
 sg13g2_xnor2_1 _4212_ (.Y(_1181_),
    .A(_1110_),
    .B(_1129_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4213_ (.Y(_1182_),
    .B1(net567),
    .B2(_1181_),
    .A2(_1131_),
    .A1(_2290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4214_ (.VDD(VPWR),
    .Y(_1183_),
    .A(_1182_),
    .VSS(VGND));
 sg13g2_o21ai_1 _4215_ (.B1(net805),
    .VDD(VPWR),
    .Y(_1184_),
    .VSS(VGND),
    .A1(net1079),
    .A2(net635));
 sg13g2_a21oi_1 _4216_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net634),
    .A2(_1183_),
    .Y(_0279_),
    .B1(net1080));
 sg13g2_nor2_1 _4217_ (.A(net779),
    .B(_2152_),
    .Y(_1185_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4218_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net779),
    .A2(\falu_i.falutop.div_inst.a[0] ),
    .Y(_1186_),
    .B1(_1185_));
 sg13g2_nor2_1 _4219_ (.A(net399),
    .B(net606),
    .Y(_1187_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4220_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net606),
    .A2(_1186_),
    .Y(_0280_),
    .B1(_1187_));
 sg13g2_nor2_1 _4221_ (.A(net780),
    .B(_2151_),
    .Y(_1188_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4222_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net780),
    .A2(net388),
    .Y(_1189_),
    .B1(_1188_));
 sg13g2_nor2_1 _4223_ (.A(net411),
    .B(net605),
    .Y(_1190_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4224_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net605),
    .A2(_1189_),
    .Y(_0281_),
    .B1(_1190_));
 sg13g2_nor2_1 _4225_ (.A(net780),
    .B(_2150_),
    .Y(_1191_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4226_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net780),
    .A2(\falu_i.falutop.div_inst.a[2] ),
    .Y(_1192_),
    .B1(_1191_));
 sg13g2_nor2_1 _4227_ (.A(net435),
    .B(net605),
    .Y(_1193_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4228_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net605),
    .A2(_1192_),
    .Y(_0282_),
    .B1(_1193_));
 sg13g2_nor2_1 _4229_ (.A(net781),
    .B(_2149_),
    .Y(_1194_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4230_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net781),
    .A2(\falu_i.falutop.div_inst.a[3] ),
    .Y(_1195_),
    .B1(_1194_));
 sg13g2_nor2_1 _4231_ (.A(net405),
    .B(net605),
    .Y(_1196_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4232_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1106_),
    .A2(_1195_),
    .Y(_0283_),
    .B1(_1196_));
 sg13g2_nor2_1 _4233_ (.A(net781),
    .B(_2148_),
    .Y(_1197_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4234_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net781),
    .A2(\falu_i.falutop.div_inst.a[4] ),
    .Y(_1198_),
    .B1(_1197_));
 sg13g2_nor2_1 _4235_ (.A(net432),
    .B(net605),
    .Y(_1199_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4236_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net606),
    .A2(_1198_),
    .Y(_0284_),
    .B1(_1199_));
 sg13g2_nor2_1 _4237_ (.A(net780),
    .B(_2147_),
    .Y(_1200_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4238_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net780),
    .A2(net465),
    .Y(_1201_),
    .B1(_1200_));
 sg13g2_nor2_1 _4239_ (.A(net542),
    .B(net605),
    .Y(_1202_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4240_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net605),
    .A2(_1201_),
    .Y(_0285_),
    .B1(_1202_));
 sg13g2_nor2_1 _4241_ (.A(net780),
    .B(_2146_),
    .Y(_1203_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4242_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net780),
    .A2(\falu_i.falutop.div_inst.a[6] ),
    .Y(_1204_),
    .B1(_1203_));
 sg13g2_nor2_1 _4243_ (.A(net396),
    .B(net606),
    .Y(_1205_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4244_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net606),
    .A2(_1204_),
    .Y(_0286_),
    .B1(_1205_));
 sg13g2_nand2_1 _4245_ (.Y(_1206_),
    .A(net498),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4246_ (.B1(_1206_),
    .VDD(VPWR),
    .Y(_0287_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1155_));
 sg13g2_nand2_1 _4247_ (.Y(_1207_),
    .A(net489),
    .B(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4248_ (.B1(_1207_),
    .VDD(VPWR),
    .Y(_0288_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1159_));
 sg13g2_nand2_1 _4249_ (.Y(_1208_),
    .A(net494),
    .B(_1105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4250_ (.B1(_1208_),
    .VDD(VPWR),
    .Y(_0289_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1163_));
 sg13g2_nand2_1 _4251_ (.Y(_1209_),
    .A(net856),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4252_ (.B1(_1209_),
    .VDD(VPWR),
    .Y(_0290_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1167_));
 sg13g2_nand2_1 _4253_ (.Y(_1210_),
    .A(net549),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4254_ (.B1(_1210_),
    .VDD(VPWR),
    .Y(_0291_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1171_));
 sg13g2_nand2_1 _4255_ (.Y(_1211_),
    .A(net931),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4256_ (.B1(_1211_),
    .VDD(VPWR),
    .Y(_0292_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1175_));
 sg13g2_nand2_1 _4257_ (.Y(_1212_),
    .A(net485),
    .B(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4258_ (.B1(_1212_),
    .VDD(VPWR),
    .Y(_0293_),
    .VSS(VGND),
    .A1(_1098_),
    .A2(_1179_));
 sg13g2_a22oi_1 _4259_ (.Y(_1213_),
    .B1(_1182_),
    .B2(_1097_),
    .A2(net607),
    .A1(net879),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4260_ (.VDD(VPWR),
    .Y(_0294_),
    .A(net880),
    .VSS(VGND));
 sg13g2_nor2_2 _4261_ (.A(_2296_),
    .B(_2305_),
    .Y(_1214_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4262_ (.Y(_1215_),
    .A(net724),
    .B(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4263_ (.A(net722),
    .B(net750),
    .Y(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4264_ (.A(_1214_),
    .B(_1216_),
    .Y(_1217_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4265_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1218_),
    .B(_1216_),
    .A(_1214_));
 sg13g2_and2_1 _4266_ (.A(net744),
    .B(net770),
    .X(_1219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4267_ (.Y(_1220_),
    .A(net745),
    .B(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4268_ (.A(net744),
    .B(net770),
    .Y(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4269_ (.A(_1219_),
    .B(_1221_),
    .Y(_1222_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4270_ (.VDD(VPWR),
    .Y(_1223_),
    .A(_1222_),
    .VSS(VGND));
 sg13g2_and2_1 _4271_ (.A(net732),
    .B(net757),
    .X(_1224_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4272_ (.B(net760),
    .A(net730),
    .X(_1225_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4273_ (.A(net739),
    .B(net764),
    .Y(_1226_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4274_ (.A(net737),
    .B(net763),
    .X(_1227_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4275_ (.Y(_1228_),
    .A(net736),
    .B(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4276_ (.A(_1226_),
    .B(_1227_),
    .Y(_1229_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4277_ (.Y(_1230_),
    .B(_1228_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1226_));
 sg13g2_nor2_2 _4278_ (.A(\falu_i.falutop.alu_data_in[9] ),
    .B(net767),
    .Y(_1231_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4279_ (.A(net707),
    .B(_2304_),
    .Y(_1232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4280_ (.Y(_1233_),
    .A(net741),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4281_ (.A(_1231_),
    .B(_1232_),
    .Y(_1234_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4282_ (.Y(_1235_),
    .B(_1233_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1231_));
 sg13g2_and2_1 _4283_ (.A(net729),
    .B(net754),
    .X(_1236_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4284_ (.Y(_1237_),
    .A(net729),
    .B(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4285_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1238_),
    .B(net754),
    .A(net729));
 sg13g2_and2_1 _4286_ (.A(_1237_),
    .B(_1238_),
    .X(_1239_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4287_ (.A(net714),
    .B(\falu_i.falutop.alu_data_in[7] ),
    .Y(_1240_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4288_ (.Y(_1241_),
    .A(net714),
    .B(\falu_i.falutop.alu_data_in[7] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4289_ (.Y(_1242_),
    .B(_1241_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1240_));
 sg13g2_and2_1 _4290_ (.A(net717),
    .B(net747),
    .X(_1243_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4291_ (.Y(_1244_),
    .A(net720),
    .B(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4292_ (.A(net717),
    .B(net747),
    .Y(_1245_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4293_ (.A(_1243_),
    .B(_1245_),
    .Y(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4294_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1247_),
    .B(_1245_),
    .A(_1243_));
 sg13g2_xnor2_1 _4295_ (.Y(_1248_),
    .A(net632),
    .B(_1246_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4296_ (.Y(_1249_),
    .A(_1239_),
    .B(_1248_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4297_ (.B(_1248_),
    .A(_1239_),
    .X(_1250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4298_ (.A(_1234_),
    .B(_1250_),
    .X(_1251_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4299_ (.Y(_1252_),
    .A(_1235_),
    .B(_1250_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4300_ (.Y(_1253_),
    .A(_1230_),
    .B(_1252_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4301_ (.A(_1225_),
    .B(_1253_),
    .X(_1254_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4302_ (.B(_1253_),
    .A(_1225_),
    .X(_1255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4303_ (.Y(_1256_),
    .A(_1222_),
    .B(_1255_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4304_ (.Y(_1257_),
    .A(_1218_),
    .B(_1256_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4305_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1258_),
    .B(_1256_),
    .A(_1218_));
 sg13g2_nand2_2 _4306_ (.Y(_1259_),
    .A(net772),
    .B(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4307_ (.Y(_1260_),
    .A(\falu_i.falutop.alu_inst.op[1] ),
    .B(net877),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4308_ (.A(_1259_),
    .B(_1260_),
    .Y(_1261_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4309_ (.B(_1258_),
    .C(_1261_),
    .A(_1257_),
    .Y(_1262_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4310_ (.Y(_1263_),
    .B(net759),
    .A_N(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4311_ (.Y(_1264_),
    .B(net764),
    .A_N(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4312_ (.A(net740),
    .B(_2304_),
    .Y(_1265_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4313_ (.Y(_1266_),
    .A(net745),
    .B(_2301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4314_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1235_),
    .A2(_1266_),
    .Y(_1267_),
    .B1(_1265_));
 sg13g2_or2_1 _4315_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1268_),
    .B(_1267_),
    .A(_1229_));
 sg13g2_a21o_1 _4316_ (.A2(_1268_),
    .A1(_1264_),
    .B1(_1225_),
    .X(_1269_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4317_ (.A2(_1269_),
    .A1(_1263_),
    .B1(_1239_),
    .X(_1270_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4318_ (.Y(_1271_),
    .B(net752),
    .A_N(net729),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4319_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1270_),
    .A2(_1271_),
    .Y(_1272_),
    .B1(_1217_));
 sg13g2_a21oi_1 _4320_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2296_),
    .A2(net750),
    .Y(_1273_),
    .B1(_1272_));
 sg13g2_and3_1 _4321_ (.X(_1274_),
    .A(net632),
    .B(_1247_),
    .C(_1273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4322_ (.A(net714),
    .B(net705),
    .Y(_1275_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4323_ (.A(\falu_i.falutop.alu_data_in[7] ),
    .B_N(net714),
    .Y(_1276_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4324_ (.A(_2297_),
    .B(net747),
    .C(_1275_),
    .Y(_1277_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4325_ (.A(_1274_),
    .B(_1276_),
    .C(_1277_),
    .Y(_1278_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4326_ (.Y(_1279_),
    .A(\falu_i.falutop.alu_inst.op[1] ),
    .B(_2298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4327_ (.A(net772),
    .B(_1279_),
    .Y(_1280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _4328_ (.A(net772),
    .B(_2300_),
    .C(_1279_),
    .Y(_1281_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4329_ (.Y(_1282_),
    .A(\falu_i.falutop.alu_inst.op[3] ),
    .B(_1280_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4330_ (.A0(net770),
    .A1(net744),
    .S(net566),
    .X(_1283_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4331_ (.A(net716),
    .B(net710),
    .Y(_1284_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4332_ (.A(net730),
    .B(net736),
    .Y(_1285_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4333_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1286_),
    .B(net725),
    .A(net721));
 sg13g2_nor2_1 _4334_ (.A(_1285_),
    .B(_1286_),
    .Y(_1287_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _4335_ (.A(_1287_),
    .B_N(_1284_),
    .Y(_1288_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _4336_ (.A(net716),
    .B(net710),
    .C(_1286_),
    .Y(_1289_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4337_ (.A(net707),
    .B(net735),
    .Y(_1290_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4338_ (.B1(_1289_),
    .VDD(VPWR),
    .Y(_1291_),
    .VSS(VGND),
    .A1(net730),
    .A2(_1290_));
 sg13g2_nand2b_1 _4339_ (.Y(_1292_),
    .B(_1291_),
    .A_N(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4340_ (.A(_2296_),
    .B(net716),
    .Y(_1293_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4341_ (.Y(_1294_),
    .B(_2296_),
    .A_N(_1292_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4342_ (.A(_1292_),
    .B(_1293_),
    .Y(_1295_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4343_ (.Y(_1296_),
    .A(net743),
    .B(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4344_ (.B1(_1296_),
    .VDD(VPWR),
    .Y(_1297_),
    .VSS(VGND),
    .A1(net707),
    .A2(net587));
 sg13g2_nand4_1 _4345_ (.B(\falu_i.falutop.alu_inst.op[0] ),
    .C(_2299_),
    .A(\falu_i.falutop.alu_inst.op[1] ),
    .Y(_1298_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net771));
 sg13g2_nor2_2 _4346_ (.A(_1289_),
    .B(_1298_),
    .Y(_1299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4347_ (.A0(net730),
    .A1(net735),
    .S(net587),
    .X(_1300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4348_ (.A0(_1300_),
    .A1(_1297_),
    .S(_1288_),
    .X(_1301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4349_ (.A(\falu_i.falutop.alu_inst.op[1] ),
    .B(\falu_i.falutop.alu_inst.op[0] ),
    .Y(_1302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _4350_ (.A(\falu_i.falutop.alu_inst.op[1] ),
    .B(\falu_i.falutop.alu_inst.op[0] ),
    .C(net771),
    .Y(_1303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4351_ (.Y(_1304_),
    .B(\falu_i.falutop.alu_inst.op[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(\falu_i.falutop.alu_inst.op[1] ));
 sg13g2_nor2_1 _4352_ (.A(net772),
    .B(net771),
    .Y(_1305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_2 _4353_ (.A(_1304_),
    .B_N(_1305_),
    .Y(_1306_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4354_ (.B1(_1220_),
    .VDD(VPWR),
    .Y(_1307_),
    .VSS(VGND),
    .A1(_1303_),
    .A2(net631));
 sg13g2_nand2_1 _4355_ (.Y(_1308_),
    .A(net726),
    .B(_1219_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _4356_ (.A(net772),
    .B(_2300_),
    .C(_1304_),
    .Y(_1309_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4357_ (.VDD(VPWR),
    .Y(_1310_),
    .A(_1309_),
    .VSS(VGND));
 sg13g2_or2_1 _4358_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1311_),
    .B(net770),
    .A(net726));
 sg13g2_nand3_1 _4359_ (.B(_1309_),
    .C(_1311_),
    .A(_1308_),
    .Y(_1312_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4360_ (.A(_1260_),
    .B_N(_1305_),
    .Y(_1313_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_2 _4361_ (.Y(_1314_),
    .B(_1305_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1260_));
 sg13g2_nand3_1 _4362_ (.B(_1312_),
    .C(_1314_),
    .A(_1307_),
    .Y(_1315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4363_ (.Y(_1316_),
    .B(_1315_),
    .A_N(_1221_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4364_ (.A(_1259_),
    .B(_1279_),
    .Y(_1317_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4365_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1318_),
    .B(_1279_),
    .A(_1259_));
 sg13g2_nor3_2 _4366_ (.A(net772),
    .B(net771),
    .C(_1279_),
    .Y(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4367_ (.B1(_1219_),
    .VDD(VPWR),
    .Y(_1320_),
    .VSS(VGND),
    .A1(net615),
    .A2(_1319_));
 sg13g2_nand2_2 _4368_ (.Y(_1321_),
    .A(\falu_i.falutop.alu_inst.op[2] ),
    .B(_2300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4369_ (.A(_1260_),
    .B(_1321_),
    .Y(_1322_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4370_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1323_),
    .B(_1321_),
    .A(_1260_));
 sg13g2_nor2_2 _4371_ (.A(_1279_),
    .B(_1321_),
    .Y(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4372_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1325_),
    .B(_1321_),
    .A(_1279_));
 sg13g2_o21ai_1 _4373_ (.B1(_1323_),
    .VDD(VPWR),
    .Y(_1326_),
    .VSS(VGND),
    .A1(net744),
    .A2(_1325_));
 sg13g2_nor2_2 _4374_ (.A(_1304_),
    .B(_1321_),
    .Y(_1327_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4375_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1220_),
    .C1(net640),
    .B1(_1327_),
    .A1(_1223_),
    .Y(_1328_),
    .A2(_1326_));
 sg13g2_nor2b_1 _4376_ (.A(_1259_),
    .B_N(_1302_),
    .Y(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4377_ (.Y(_1330_),
    .B(net730),
    .A_N(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4378_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net707),
    .A2(_1330_),
    .Y(_1331_),
    .B1(net743));
 sg13g2_nor2_1 _4379_ (.A(net743),
    .B(net740),
    .Y(_1332_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4380_ (.A(_1285_),
    .B(_1332_),
    .X(_1333_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4381_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2297_),
    .A2(net710),
    .Y(_1334_),
    .B1(net722));
 sg13g2_nor2_1 _4382_ (.A(net726),
    .B(_1334_),
    .Y(_1335_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4383_ (.A2(_1335_),
    .A1(_1333_),
    .B1(_1331_),
    .X(_1336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4384_ (.B(net771),
    .C(_1302_),
    .A(_2299_),
    .Y(_1337_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4385_ (.VDD(VPWR),
    .Y(_1338_),
    .A(_1337_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4386_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net743),
    .A2(net707),
    .Y(_1339_),
    .B1(net735));
 sg13g2_nand2b_1 _4387_ (.Y(_1340_),
    .B(_1289_),
    .A_N(_1339_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4388_ (.A(net710),
    .B(_1293_),
    .Y(_1341_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4389_ (.B1(_1341_),
    .VDD(VPWR),
    .Y(_1342_),
    .VSS(VGND),
    .A1(net725),
    .A2(net717));
 sg13g2_o21ai_1 _4390_ (.B1(_1342_),
    .VDD(VPWR),
    .Y(_1343_),
    .VSS(VGND),
    .A1(net731),
    .A2(_1340_));
 sg13g2_a22oi_1 _4391_ (.Y(_1344_),
    .B1(_1338_),
    .B2(_1343_),
    .A2(_1336_),
    .A1(_1329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4392_ (.B(_1320_),
    .C(_1328_),
    .A(_1316_),
    .Y(_1345_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1344_));
 sg13g2_a221oi_1 _4393_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1301_),
    .C1(_1345_),
    .B1(_1299_),
    .A1(net616),
    .Y(_1346_),
    .A2(_1283_));
 sg13g2_nand2_1 _4394_ (.Y(_1347_),
    .A(_1262_),
    .B(_1346_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4395_ (.B1(_1347_),
    .VDD(VPWR),
    .Y(_1348_),
    .VSS(VGND),
    .A1(\falu_i.falutop.div_inst.val[0] ),
    .A2(_1074_));
 sg13g2_o21ai_1 _4396_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1349_),
    .VSS(VGND),
    .A1(net1022),
    .A2(net628));
 sg13g2_a21oi_1 _4397_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net628),
    .A2(_1348_),
    .Y(_0295_),
    .B1(_1349_));
 sg13g2_o21ai_1 _4398_ (.B1(_1249_),
    .VDD(VPWR),
    .Y(_1350_),
    .VSS(VGND),
    .A1(net632),
    .A2(_1247_));
 sg13g2_a21oi_1 _4399_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1229_),
    .A2(_1252_),
    .Y(_1351_),
    .B1(_1251_));
 sg13g2_inv_1 _4400_ (.VDD(VPWR),
    .Y(_1352_),
    .A(_1351_),
    .VSS(VGND));
 sg13g2_nand2_1 _4401_ (.Y(_1353_),
    .A(_1350_),
    .B(_1352_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4402_ (.Y(_1354_),
    .A(_1350_),
    .B(_1351_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4403_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1222_),
    .A2(_1255_),
    .Y(_1355_),
    .B1(_1254_));
 sg13g2_nand2b_1 _4404_ (.Y(_1356_),
    .B(_1354_),
    .A_N(_1355_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4405_ (.B(_1355_),
    .A(_1354_),
    .X(_1357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4406_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1358_),
    .B(_1357_),
    .A(_1258_));
 sg13g2_nand2_1 _4407_ (.Y(_1359_),
    .A(_1258_),
    .B(_1357_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4408_ (.B(_1358_),
    .C(_1359_),
    .A(_1261_),
    .Y(_1360_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4409_ (.B1(net616),
    .VDD(VPWR),
    .Y(_1361_),
    .VSS(VGND),
    .A1(net767),
    .A2(net566));
 sg13g2_a21oi_1 _4410_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net707),
    .A2(net566),
    .Y(_1362_),
    .B1(_1361_));
 sg13g2_nor2_2 _4411_ (.A(_1288_),
    .B(_1298_),
    .Y(_1363_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _4412_ (.B(_1363_),
    .C(net743),
    .Y(_1364_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(net587));
 sg13g2_nand2b_1 _4413_ (.Y(_1365_),
    .B(_1364_),
    .A_N(_1299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4414_ (.A0(net725),
    .A1(net730),
    .S(net587),
    .X(_1366_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4415_ (.A(net736),
    .B(net587),
    .Y(_1367_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4416_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net707),
    .A2(net587),
    .Y(_1368_),
    .B1(_1367_));
 sg13g2_mux2_1 _4417_ (.A0(_1366_),
    .A1(_1368_),
    .S(_1284_),
    .X(_1369_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4418_ (.B1(_1365_),
    .VDD(VPWR),
    .Y(_1370_),
    .VSS(VGND),
    .A1(_1289_),
    .A2(_1369_));
 sg13g2_nand2b_1 _4419_ (.Y(_1371_),
    .B(_1332_),
    .A_N(_1286_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4420_ (.X(_1372_),
    .A(_1288_),
    .B(_1338_),
    .C(_1371_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4421_ (.A(_2299_),
    .B(_1303_),
    .X(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4422_ (.Y(_1374_),
    .A(_2299_),
    .B(_1303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4423_ (.Y(_1375_),
    .A(_1219_),
    .B(_1235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4424_ (.B1(_1285_),
    .VDD(VPWR),
    .Y(_1376_),
    .VSS(VGND),
    .A1(_1284_),
    .A2(_1286_));
 sg13g2_and3_1 _4425_ (.X(_1377_),
    .A(_1329_),
    .B(_1332_),
    .C(_1376_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4426_ (.A(_1220_),
    .B(_1233_),
    .Y(_1378_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4427_ (.VDD(VPWR),
    .Y(_1379_),
    .A(_1378_),
    .VSS(VGND));
 sg13g2_a22oi_1 _4428_ (.Y(_1380_),
    .B1(net766),
    .B2(net745),
    .A2(net769),
    .A1(net741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4429_ (.A(_1318_),
    .B(_1378_),
    .C(_1380_),
    .Y(_1381_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4430_ (.Y(_1382_),
    .B1(_1324_),
    .B2(_1231_),
    .A2(_1322_),
    .A1(_1235_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4431_ (.A(net772),
    .B(_1303_),
    .X(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4432_ (.Y(_1384_),
    .A(_1234_),
    .B(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4433_ (.B(_1266_),
    .A(_1235_),
    .X(_1385_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4434_ (.B1(_1384_),
    .VDD(VPWR),
    .Y(_1386_),
    .VSS(VGND),
    .A1(_1231_),
    .A2(_1314_));
 sg13g2_a22oi_1 _4435_ (.Y(_1387_),
    .B1(_1385_),
    .B2(net631),
    .A2(_1375_),
    .A1(_1373_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4436_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1233_),
    .A2(_1327_),
    .Y(_1388_),
    .B1(net640));
 sg13g2_a21oi_1 _4437_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1232_),
    .A2(_1319_),
    .Y(_1389_),
    .B1(_1381_));
 sg13g2_nand4_1 _4438_ (.B(_1387_),
    .C(_1388_),
    .A(_1382_),
    .Y(_1390_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1389_));
 sg13g2_nor4_1 _4439_ (.A(_1372_),
    .B(_1377_),
    .C(_1386_),
    .D(_1390_),
    .Y(_1391_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4440_ (.Y(_1392_),
    .A(net728),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4441_ (.Y(_1393_),
    .A(net726),
    .B(_1232_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4442_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net740),
    .A2(net726),
    .Y(_1394_),
    .B1(net767));
 sg13g2_nand2b_1 _4443_ (.Y(_1395_),
    .B(_1393_),
    .A_N(_1394_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4444_ (.Y(_1396_),
    .A(net744),
    .B(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4445_ (.A(_1395_),
    .B(_1396_),
    .Y(_1397_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4446_ (.Y(_1398_),
    .A(_1395_),
    .B(_1396_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4447_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1399_),
    .B(_1398_),
    .A(_1308_));
 sg13g2_a21oi_1 _4448_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1308_),
    .A2(_1398_),
    .Y(_1400_),
    .B1(_1310_));
 sg13g2_a21oi_1 _4449_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1399_),
    .A2(_1400_),
    .Y(_1401_),
    .B1(_1362_));
 sg13g2_nand4_1 _4450_ (.B(_1370_),
    .C(_1391_),
    .A(_1360_),
    .Y(_1402_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1401_));
 sg13g2_o21ai_1 _4451_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1403_),
    .VSS(VGND),
    .A1(net1057),
    .A2(net628));
 sg13g2_xor2_1 _4452_ (.B(net776),
    .A(\falu_i.falutop.data_in[7] ),
    .X(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4453_ (.Y(_1405_),
    .A(\falu_i.falutop.div_inst.val[0] ),
    .B(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4454_ (.Y(_1406_),
    .A(net380),
    .B(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4455_ (.Y(_1407_),
    .A(net939),
    .B(_1405_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4456_ (.B1(_1402_),
    .VDD(VPWR),
    .Y(_1408_),
    .VSS(VGND),
    .A1(_1406_),
    .A2(_1407_));
 sg13g2_nor2_1 _4457_ (.A(_1403_),
    .B(_1408_),
    .Y(_0296_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4458_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1409_),
    .B(_1358_),
    .A(_1353_));
 sg13g2_inv_1 _4459_ (.VDD(VPWR),
    .Y(_1410_),
    .A(_1409_),
    .VSS(VGND));
 sg13g2_nand3_1 _4460_ (.B(_1356_),
    .C(_1358_),
    .A(_1353_),
    .Y(_1411_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4461_ (.B(_1409_),
    .C(_1411_),
    .A(_1261_),
    .Y(_1412_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4462_ (.A0(net765),
    .A1(net736),
    .S(net566),
    .X(_1413_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4463_ (.Y(_1414_),
    .A(net743),
    .B(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4464_ (.B(net725),
    .C(net765),
    .A(net735),
    .Y(_1415_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4465_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net735),
    .A2(net725),
    .Y(_1416_),
    .B1(net765));
 sg13g2_nor2b_1 _4466_ (.A(_1416_),
    .B_N(_1415_),
    .Y(_1417_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4467_ (.Y(_1418_),
    .A(net740),
    .B(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4468_ (.B(_1418_),
    .A(_1417_),
    .X(_1419_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4469_ (.B(_1419_),
    .A(_1393_),
    .X(_1420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4470_ (.Y(_1421_),
    .B(_1420_),
    .A_N(_1414_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4471_ (.Y(_1422_),
    .A(_1414_),
    .B(_1420_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4472_ (.Y(_1423_),
    .A(_1397_),
    .B(_1422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4473_ (.Y(_1424_),
    .A(_1397_),
    .B(_1422_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4474_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1425_),
    .B(_1424_),
    .A(_1399_));
 sg13g2_a21oi_1 _4475_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1399_),
    .A2(_1424_),
    .Y(_1426_),
    .B1(_1310_));
 sg13g2_a21oi_1 _4476_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1219_),
    .A2(_1234_),
    .Y(_1427_),
    .B1(_1232_));
 sg13g2_nand2_1 _4477_ (.Y(_1428_),
    .A(net745),
    .B(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4478_ (.A(_1233_),
    .B(_1428_),
    .Y(_1429_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4479_ (.B(_1428_),
    .A(_1233_),
    .X(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4480_ (.X(_1431_),
    .A(net737),
    .B(net769),
    .C(_1430_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4481_ (.VDD(VPWR),
    .Y(_1432_),
    .A(_1431_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4482_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net737),
    .A2(net769),
    .Y(_1433_),
    .B1(_1430_));
 sg13g2_nor3_1 _4483_ (.A(_1379_),
    .B(_1431_),
    .C(_1433_),
    .Y(_1434_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4484_ (.B1(_1379_),
    .VDD(VPWR),
    .Y(_1435_),
    .VSS(VGND),
    .A1(_1431_),
    .A2(_1433_));
 sg13g2_nand2_1 _4485_ (.Y(_1436_),
    .A(net615),
    .B(_1435_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4486_ (.A(_1434_),
    .B(_1436_),
    .Y(_1437_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4487_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1291_),
    .A2(_1340_),
    .Y(_1438_),
    .B1(_1337_));
 sg13g2_nand3b_1 _4488_ (.B(_1329_),
    .C(_1333_),
    .Y(_1439_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1289_));
 sg13g2_nand2_1 _4489_ (.Y(_1440_),
    .A(_1229_),
    .B(_1267_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4490_ (.B(net631),
    .C(_1440_),
    .A(_1268_),
    .Y(_1441_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4491_ (.B1(_1228_),
    .VDD(VPWR),
    .Y(_1442_),
    .VSS(VGND),
    .A1(_1304_),
    .A2(_1321_));
 sg13g2_o21ai_1 _4492_ (.B1(_1442_),
    .VDD(VPWR),
    .Y(_1443_),
    .VSS(VGND),
    .A1(_1228_),
    .A2(_1319_));
 sg13g2_xnor2_1 _4493_ (.Y(_1444_),
    .A(_1230_),
    .B(_1427_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4494_ (.Y(_1445_),
    .A(_1229_),
    .B(_1383_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4495_ (.B1(_1441_),
    .VDD(VPWR),
    .Y(_1446_),
    .VSS(VGND),
    .A1(_1374_),
    .A2(_1444_));
 sg13g2_o21ai_1 _4496_ (.B1(_1074_),
    .VDD(VPWR),
    .Y(_1447_),
    .VSS(VGND),
    .A1(_1226_),
    .A2(_1314_));
 sg13g2_a221oi_1 _4497_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1226_),
    .C1(_1447_),
    .B1(_1324_),
    .A1(_1230_),
    .Y(_1448_),
    .A2(_1322_));
 sg13g2_nand4_1 _4498_ (.B(_1443_),
    .C(_1445_),
    .A(_1439_),
    .Y(_1449_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1448_));
 sg13g2_nor4_1 _4499_ (.A(_1437_),
    .B(_1438_),
    .C(_1446_),
    .D(_1449_),
    .Y(_1450_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4500_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1297_),
    .A2(_1363_),
    .Y(_1451_),
    .B1(_1299_));
 sg13g2_nand2b_1 _4501_ (.Y(_1452_),
    .B(net587),
    .A_N(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4502_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2296_),
    .A2(_1292_),
    .Y(_1453_),
    .B1(_1288_));
 sg13g2_a221oi_1 _4503_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1453_),
    .C1(_1289_),
    .B1(_1452_),
    .A1(_1284_),
    .Y(_1454_),
    .A2(_1300_));
 sg13g2_o21ai_1 _4504_ (.B1(_1450_),
    .VDD(VPWR),
    .Y(_1455_),
    .VSS(VGND),
    .A1(_1451_),
    .A2(_1454_));
 sg13g2_a221oi_1 _4505_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1426_),
    .C1(_1455_),
    .B1(_1425_),
    .A1(net616),
    .Y(_1456_),
    .A2(_1413_));
 sg13g2_o21ai_1 _4506_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1457_),
    .VSS(VGND),
    .A1(net1047),
    .A2(net628));
 sg13g2_o21ai_1 _4507_ (.B1(_1404_),
    .VDD(VPWR),
    .Y(_1458_),
    .VSS(VGND),
    .A1(net939),
    .A2(\falu_i.falutop.div_inst.val[0] ));
 sg13g2_or2_1 _4508_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1459_),
    .B(_1458_),
    .A(net978));
 sg13g2_a21oi_1 _4509_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net978),
    .A2(_1458_),
    .Y(_1460_),
    .B1(_1406_));
 sg13g2_a221oi_1 _4510_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1460_),
    .C1(_1457_),
    .B1(_1459_),
    .A1(_1412_),
    .Y(_0297_),
    .A2(_1456_));
 sg13g2_mux2_1 _4511_ (.A0(net760),
    .A1(net730),
    .S(net566),
    .X(_1461_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4512_ (.Y(_1462_),
    .A(net731),
    .B(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4513_ (.B1(_1421_),
    .VDD(VPWR),
    .Y(_1463_),
    .VSS(VGND),
    .A1(_1393_),
    .A2(_1419_));
 sg13g2_nand2_1 _4514_ (.Y(_1464_),
    .A(net743),
    .B(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4515_ (.B1(_1415_),
    .VDD(VPWR),
    .Y(_1465_),
    .VSS(VGND),
    .A1(_1416_),
    .A2(_1418_));
 sg13g2_nand2_1 _4516_ (.Y(_1466_),
    .A(net740),
    .B(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4517_ (.A(net735),
    .B(net760),
    .X(_1467_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4518_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net735),
    .A2(net721),
    .Y(_1468_),
    .B1(net760));
 sg13g2_a21o_1 _4519_ (.A2(_1467_),
    .A1(net721),
    .B1(_1468_),
    .X(_1469_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4520_ (.A(_1466_),
    .B(_1469_),
    .Y(_1470_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4521_ (.B(_1469_),
    .A(_1466_),
    .X(_1471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4522_ (.Y(_1472_),
    .A(_1465_),
    .B(_1471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4523_ (.Y(_1473_),
    .A(_1465_),
    .B(_1471_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4524_ (.B(_1473_),
    .A(_1464_),
    .X(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4525_ (.Y(_1475_),
    .A(_1463_),
    .B(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4526_ (.Y(_1476_),
    .A(_1463_),
    .B(_1474_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4527_ (.B(_1476_),
    .A(_1462_),
    .X(_1477_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4528_ (.Y(_1478_),
    .A(_1423_),
    .B(_1425_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4529_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1479_),
    .B(_1478_),
    .A(_1477_));
 sg13g2_nand2_1 _4530_ (.Y(_1480_),
    .A(_1477_),
    .B(_1478_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4531_ (.B(_1479_),
    .C(_1480_),
    .A(_1309_),
    .Y(_1481_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4532_ (.Y(_1482_),
    .A(net732),
    .B(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4533_ (.Y(_1483_),
    .A(net737),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4534_ (.A(net745),
    .B(net741),
    .C(net763),
    .D(net757),
    .X(_1484_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4535_ (.B(net741),
    .C(net762),
    .A(net745),
    .Y(_1485_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net756));
 sg13g2_a22oi_1 _4536_ (.Y(_1486_),
    .B1(net756),
    .B2(net745),
    .A2(net762),
    .A1(net741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4537_ (.A(_1483_),
    .B(_1484_),
    .C(_1486_),
    .X(_1487_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4538_ (.B1(_1483_),
    .VDD(VPWR),
    .Y(_1488_),
    .VSS(VGND),
    .A1(_1484_),
    .A2(_1486_));
 sg13g2_and3_1 _4539_ (.X(_1489_),
    .A(_1429_),
    .B(_1487_),
    .C(_1488_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4540_ (.B(_1487_),
    .C(_1488_),
    .A(_1429_),
    .Y(_1490_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4541_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1487_),
    .A2(_1488_),
    .Y(_1491_),
    .B1(_1429_));
 sg13g2_nor2_1 _4542_ (.A(_1489_),
    .B(_1491_),
    .Y(_1492_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4543_ (.B(_1492_),
    .A(_1482_),
    .X(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4544_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1494_),
    .B(_1493_),
    .A(_1432_));
 sg13g2_xnor2_1 _4545_ (.Y(_1495_),
    .A(_1431_),
    .B(_1493_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4546_ (.A(_1434_),
    .B(_1495_),
    .X(_1496_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4547_ (.A(_1318_),
    .B(_1496_),
    .Y(_1497_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4548_ (.B1(_1497_),
    .VDD(VPWR),
    .Y(_1498_),
    .VSS(VGND),
    .A1(_1434_),
    .A2(_1495_));
 sg13g2_a221oi_1 _4549_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1288_),
    .C1(_1289_),
    .B1(_1366_),
    .A1(net716),
    .Y(_1499_),
    .A2(_1294_));
 sg13g2_nor2_1 _4550_ (.A(_1295_),
    .B(_1298_),
    .Y(_1500_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4551_ (.B(_1288_),
    .C(_1500_),
    .A(net744),
    .Y(_1501_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4552_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1363_),
    .A2(_1368_),
    .Y(_1502_),
    .B1(_1299_));
 sg13g2_a21o_1 _4553_ (.A2(_1502_),
    .A1(_1501_),
    .B1(_1499_),
    .X(_1503_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4554_ (.B(_1264_),
    .C(_1268_),
    .A(_1225_),
    .Y(_1504_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4555_ (.A(_1269_),
    .B(_1504_),
    .X(_1505_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4556_ (.B1(_1228_),
    .VDD(VPWR),
    .Y(_1506_),
    .VSS(VGND),
    .A1(_1230_),
    .A2(_1427_));
 sg13g2_and2_1 _4557_ (.A(_1225_),
    .B(_1506_),
    .X(_1507_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4558_ (.B(_1506_),
    .A(_1225_),
    .X(_1508_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4559_ (.B1(_1314_),
    .VDD(VPWR),
    .Y(_1509_),
    .VSS(VGND),
    .A1(net734),
    .A2(net759));
 sg13g2_or3_1 _4560_ (.A(net734),
    .B(net759),
    .C(_1324_),
    .X(_1510_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4561_ (.A(_1225_),
    .B(_1323_),
    .Y(_1511_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4562_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1510_),
    .C1(_1511_),
    .B1(_1509_),
    .A1(_1225_),
    .Y(_1512_),
    .A2(_1383_));
 sg13g2_nand4_1 _4563_ (.B(_1289_),
    .C(_1302_),
    .A(net771),
    .Y(_1513_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1333_));
 sg13g2_nand2_1 _4564_ (.Y(_1514_),
    .A(_1224_),
    .B(_1319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4565_ (.A(_1224_),
    .B(_1304_),
    .C(_1321_),
    .Y(_1515_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4566_ (.A(net640),
    .B(_1515_),
    .Y(_1516_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4567_ (.B(_1513_),
    .C(_1514_),
    .A(_1512_),
    .Y(_1517_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1516_));
 sg13g2_a221oi_1 _4568_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1373_),
    .C1(_1517_),
    .B1(_1508_),
    .A1(net631),
    .Y(_1518_),
    .A2(_1505_));
 sg13g2_nand4_1 _4569_ (.B(_1498_),
    .C(_1503_),
    .A(_1481_),
    .Y(_1519_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1518_));
 sg13g2_a221oi_1 _4570_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net616),
    .C1(_1519_),
    .B1(_1461_),
    .A1(_1261_),
    .Y(_1520_),
    .A2(_1410_));
 sg13g2_o21ai_1 _4571_ (.B1(net819),
    .VDD(VPWR),
    .Y(_1521_),
    .VSS(VGND),
    .A1(net1089),
    .A2(net629));
 sg13g2_nand2_1 _4572_ (.Y(_1522_),
    .A(\falu_i.falutop.div_inst.val[2] ),
    .B(_1404_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4573_ (.A(_1458_),
    .B(_1522_),
    .X(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4574_ (.Y(_1524_),
    .B(net947),
    .A_N(_1523_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4575_ (.Y(_1525_),
    .B(_1523_),
    .A_N(net947),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4576_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1524_),
    .A2(_1525_),
    .Y(_1526_),
    .B1(_1406_));
 sg13g2_nor3_1 _4577_ (.A(_1520_),
    .B(_1521_),
    .C(_1526_),
    .Y(_0298_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4578_ (.Y(_1527_),
    .A(net731),
    .B(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4579_ (.Y(_1528_),
    .A(net740),
    .B(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4580_ (.Y(_1529_),
    .A(net737),
    .B(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4581_ (.B(net717),
    .C(net754),
    .A(net736),
    .Y(_1530_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4582_ (.A2(net717),
    .A1(net736),
    .B1(net754),
    .X(_1531_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4583_ (.A(_1530_),
    .B(_1531_),
    .X(_1532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4584_ (.Y(_1533_),
    .B(_1532_),
    .A_N(_1528_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4585_ (.Y(_1534_),
    .A(_1528_),
    .B(_1532_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4586_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net721),
    .A2(_1467_),
    .Y(_1535_),
    .B1(_1470_));
 sg13g2_nand2b_1 _4587_ (.Y(_1536_),
    .B(_1534_),
    .A_N(_1535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4588_ (.Y(_1537_),
    .A(_1534_),
    .B(_1535_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4589_ (.B1(_1472_),
    .VDD(VPWR),
    .Y(_1538_),
    .VSS(VGND),
    .A1(_1464_),
    .A2(_1473_));
 sg13g2_xor2_1 _4590_ (.B(_1538_),
    .A(_1537_),
    .X(_1539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4591_ (.A(_1527_),
    .B_N(_1539_),
    .Y(_1540_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4592_ (.Y(_1541_),
    .A(_1527_),
    .B(_1539_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4593_ (.B1(_1475_),
    .VDD(VPWR),
    .Y(_1542_),
    .VSS(VGND),
    .A1(_1462_),
    .A2(_1476_));
 sg13g2_and2_1 _4594_ (.A(_1541_),
    .B(_1542_),
    .X(_1543_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4595_ (.B(_1542_),
    .A(_1541_),
    .X(_1544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4596_ (.A(_1480_),
    .B_N(_1544_),
    .Y(_1545_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4597_ (.Y(_1546_),
    .A(_1480_),
    .B(_1544_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _4598_ (.A0(net754),
    .A1(net726),
    .S(net566),
    .X(_1547_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4599_ (.B1(_1490_),
    .VDD(VPWR),
    .Y(_1548_),
    .VSS(VGND),
    .A1(_1482_),
    .A2(_1491_));
 sg13g2_nor2_2 _4600_ (.A(_1220_),
    .B(_1237_),
    .Y(_1549_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4601_ (.VDD(VPWR),
    .Y(_1550_),
    .A(_1549_),
    .VSS(VGND));
 sg13g2_a22oi_1 _4602_ (.Y(_1551_),
    .B1(net752),
    .B2(net745),
    .A2(net770),
    .A1(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4603_ (.A(_1549_),
    .B(_1551_),
    .Y(_1552_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4604_ (.B1(_1485_),
    .VDD(VPWR),
    .Y(_1553_),
    .VSS(VGND),
    .A1(_1483_),
    .A2(_1486_));
 sg13g2_nand2_1 _4605_ (.Y(_1554_),
    .A(net732),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4606_ (.A(net741),
    .B(net737),
    .C(net762),
    .D(net756),
    .X(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4607_ (.Y(_1556_),
    .B1(net756),
    .B2(net741),
    .A2(net762),
    .A1(net737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4608_ (.A(_1554_),
    .B(_1555_),
    .C(_1556_),
    .X(_1557_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4609_ (.B1(_1554_),
    .VDD(VPWR),
    .Y(_1558_),
    .VSS(VGND),
    .A1(_1555_),
    .A2(_1556_));
 sg13g2_and3_1 _4610_ (.X(_1559_),
    .A(_1553_),
    .B(_1557_),
    .C(_1558_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4611_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1557_),
    .A2(_1558_),
    .Y(_1560_),
    .B1(_1553_));
 sg13g2_nor2_1 _4612_ (.A(_1559_),
    .B(_1560_),
    .Y(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4613_ (.Y(_1562_),
    .A(_1552_),
    .B(_1561_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4614_ (.Y(_1563_),
    .B(_1548_),
    .A_N(_1562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4615_ (.A(_1548_),
    .B_N(_1562_),
    .Y(_1564_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4616_ (.Y(_1565_),
    .A(_1548_),
    .B(_1562_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4617_ (.Y(_1566_),
    .A(_1494_),
    .B(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4618_ (.Y(_1567_),
    .A(_1496_),
    .B(_1565_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4619_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1496_),
    .A2(_1565_),
    .Y(_1568_),
    .B1(_1318_));
 sg13g2_o21ai_1 _4620_ (.B1(_1568_),
    .VDD(VPWR),
    .Y(_1569_),
    .VSS(VGND),
    .A1(_1496_),
    .A2(_1566_));
 sg13g2_nor2_1 _4621_ (.A(_1224_),
    .B(_1507_),
    .Y(_1570_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4622_ (.A(_1224_),
    .B(_1239_),
    .C(_1507_),
    .Y(_1571_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4623_ (.A(_1570_),
    .B_N(_1239_),
    .Y(_1572_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4624_ (.A(_1374_),
    .B(_1571_),
    .C(_1572_),
    .Y(_1573_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4625_ (.B1(_1074_),
    .VDD(VPWR),
    .Y(_1574_),
    .VSS(VGND),
    .A1(_1238_),
    .A2(_1325_));
 sg13g2_a22oi_1 _4626_ (.Y(_1575_),
    .B1(_1327_),
    .B2(_1237_),
    .A2(_1313_),
    .A1(_1238_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4627_ (.B1(_1575_),
    .VDD(VPWR),
    .Y(_1576_),
    .VSS(VGND),
    .A1(_1239_),
    .A2(_1323_));
 sg13g2_a221oi_1 _4628_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1239_),
    .C1(_1574_),
    .B1(_1383_),
    .A1(_1236_),
    .Y(_1577_),
    .A2(_1319_));
 sg13g2_nand2b_1 _4629_ (.Y(_1578_),
    .B(_1577_),
    .A_N(_1576_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4630_ (.A(_1500_),
    .B(_1573_),
    .C(_1578_),
    .Y(_1579_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4631_ (.B(_1263_),
    .C(_1269_),
    .A(_1239_),
    .Y(_1580_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4632_ (.B(_1306_),
    .C(_1580_),
    .A(_1270_),
    .Y(_1581_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4633_ (.B(_1579_),
    .C(_1581_),
    .A(_1569_),
    .Y(_1582_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4634_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net616),
    .C1(_1582_),
    .B1(_1547_),
    .A1(_1309_),
    .Y(_1583_),
    .A2(_1546_));
 sg13g2_o21ai_1 _4635_ (.B1(net819),
    .VDD(VPWR),
    .Y(_1584_),
    .VSS(VGND),
    .A1(net1083),
    .A2(net628));
 sg13g2_a21oi_1 _4636_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1404_),
    .A2(_1525_),
    .Y(_1585_),
    .B1(net905));
 sg13g2_nand3_1 _4637_ (.B(_1404_),
    .C(_1525_),
    .A(net905),
    .Y(_1586_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4638_ (.A(_1585_),
    .B_N(_1586_),
    .Y(_1587_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4639_ (.A(_1406_),
    .B(_1587_),
    .Y(_1588_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4640_ (.A(_1583_),
    .B(_1584_),
    .C(_1588_),
    .Y(_0299_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4641_ (.A(_1259_),
    .B(_1304_),
    .Y(_1589_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_2 _4642_ (.A(net640),
    .B(_1589_),
    .Y(_1590_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4643_ (.A(net731),
    .B(net716),
    .X(_1591_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4644_ (.X(_1592_),
    .A(net739),
    .B(net715),
    .C(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4645_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net739),
    .A2(net715),
    .Y(_1593_),
    .B1(net750));
 sg13g2_or2_1 _4646_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1594_),
    .B(_1593_),
    .A(_1592_));
 sg13g2_a21o_2 _4647_ (.A2(_1533_),
    .A1(_1530_),
    .B1(_1594_),
    .X(_1595_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4648_ (.B(_1533_),
    .C(_1594_),
    .A(_1530_),
    .Y(_1596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4649_ (.Y(_1597_),
    .A(_1595_),
    .B(_1596_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4650_ (.A(_1536_),
    .B(_1597_),
    .Y(_1598_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4651_ (.B(_1597_),
    .A(_1536_),
    .X(_1599_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4652_ (.B(_1599_),
    .A(_1591_),
    .X(_1600_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4653_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1537_),
    .A2(_1538_),
    .Y(_1601_),
    .B1(_1540_));
 sg13g2_nand2b_1 _4654_ (.Y(_1602_),
    .B(_1600_),
    .A_N(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4655_ (.Y(_1603_),
    .A(_1600_),
    .B(_1601_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4656_ (.A(_1543_),
    .B(_1545_),
    .C(_1603_),
    .Y(_1604_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4657_ (.B1(_1603_),
    .VDD(VPWR),
    .Y(_1605_),
    .VSS(VGND),
    .A1(_1543_),
    .A2(_1545_));
 sg13g2_nand2_1 _4658_ (.Y(_1606_),
    .A(_1309_),
    .B(_1605_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4659_ (.A(net750),
    .B(net565),
    .Y(_1607_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4660_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2296_),
    .A2(net565),
    .Y(_1608_),
    .B1(_1607_));
 sg13g2_nand3_1 _4661_ (.B(_1270_),
    .C(_1271_),
    .A(_1217_),
    .Y(_1609_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4662_ (.A(_1272_),
    .B_N(_1609_),
    .Y(_1610_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4663_ (.A(_1236_),
    .B(_1572_),
    .Y(_1611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4664_ (.Y(_1612_),
    .A(_1218_),
    .B(_1611_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4665_ (.A(_1216_),
    .B(_1314_),
    .Y(_1613_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4666_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1217_),
    .C1(_1363_),
    .B1(_1383_),
    .A1(_1214_),
    .Y(_1614_),
    .A2(_1319_));
 sg13g2_a22oi_1 _4667_ (.Y(_1615_),
    .B1(_1327_),
    .B2(_1215_),
    .A2(_1324_),
    .A1(_1216_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4668_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1218_),
    .A2(_1322_),
    .Y(_1616_),
    .B1(_1613_));
 sg13g2_nand3_1 _4669_ (.B(_1615_),
    .C(_1616_),
    .A(_1614_),
    .Y(_1617_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4670_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net631),
    .A2(_1610_),
    .Y(_1618_),
    .B1(_1617_));
 sg13g2_o21ai_1 _4671_ (.B1(_1618_),
    .VDD(VPWR),
    .Y(_1619_),
    .VSS(VGND),
    .A1(_1374_),
    .A2(_1612_));
 sg13g2_a21o_1 _4672_ (.A2(_1561_),
    .A1(_1552_),
    .B1(_1559_),
    .X(_1620_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4673_ (.Y(_1621_),
    .A(net746),
    .B(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4674_ (.Y(_1622_),
    .A(net724),
    .B(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4675_ (.A(_2295_),
    .B(_2301_),
    .C(_1622_),
    .Y(_1623_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4676_ (.Y(_1624_),
    .B1(net753),
    .B2(net741),
    .A2(net768),
    .A1(net723),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4677_ (.A(_1621_),
    .B(_1623_),
    .C(_1624_),
    .Y(_1625_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4678_ (.B1(_1621_),
    .VDD(VPWR),
    .Y(_1626_),
    .VSS(VGND),
    .A1(_1623_),
    .A2(_1624_));
 sg13g2_nand2b_2 _4679_ (.Y(_1627_),
    .B(_1626_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1625_));
 sg13g2_nand2b_1 _4680_ (.Y(_1628_),
    .B(_1557_),
    .A_N(_1555_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4681_ (.B(net738),
    .C(net763),
    .A(net732),
    .Y(_1629_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net756));
 sg13g2_a22oi_1 _4682_ (.Y(_1630_),
    .B1(net756),
    .B2(net737),
    .A2(net762),
    .A1(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4683_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1224_),
    .A2(_1227_),
    .Y(_1631_),
    .B1(_1630_));
 sg13g2_xor2_1 _4684_ (.B(_1631_),
    .A(_1392_),
    .X(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4685_ (.Y(_1633_),
    .B(_1628_),
    .A_N(_1632_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4686_ (.B(_1632_),
    .A(_1628_),
    .X(_1634_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4687_ (.B(_1634_),
    .A(_1627_),
    .X(_1635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4688_ (.Y(_1636_),
    .A(_1620_),
    .B(_1635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4689_ (.Y(_1637_),
    .A(_1620_),
    .B(_1635_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4690_ (.Y(_1638_),
    .A(_1549_),
    .B(_1637_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4691_ (.B1(_1563_),
    .VDD(VPWR),
    .Y(_1639_),
    .VSS(VGND),
    .A1(_1494_),
    .A2(_1564_));
 sg13g2_xnor2_1 _4692_ (.Y(_1640_),
    .A(_1638_),
    .B(_1639_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4693_ (.B(_1640_),
    .A(_1567_),
    .X(_1641_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4694_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net615),
    .C1(_1619_),
    .B1(_1641_),
    .A1(net616),
    .Y(_1642_),
    .A2(_1608_));
 sg13g2_o21ai_1 _4695_ (.B1(_1642_),
    .VDD(VPWR),
    .Y(_1643_),
    .VSS(VGND),
    .A1(_1604_),
    .A2(_1606_));
 sg13g2_nor2b_1 _4696_ (.A(_1585_),
    .B_N(_1404_),
    .Y(_1644_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4697_ (.A(net937),
    .B(_1644_),
    .Y(_1645_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4698_ (.VDD(VPWR),
    .Y(_1646_),
    .A(_1645_),
    .VSS(VGND));
 sg13g2_a21oi_1 _4699_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net937),
    .A2(_1644_),
    .Y(_1647_),
    .B1(_1074_));
 sg13g2_a221oi_1 _4700_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1647_),
    .C1(_1075_),
    .B1(_1646_),
    .A1(net614),
    .Y(_1648_),
    .A2(_1643_));
 sg13g2_o21ai_1 _4701_ (.B1(net819),
    .VDD(VPWR),
    .Y(_1649_),
    .VSS(VGND),
    .A1(net1084),
    .A2(net628));
 sg13g2_nor2_1 _4702_ (.A(_1648_),
    .B(_1649_),
    .Y(_0300_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4703_ (.B1(net819),
    .VDD(VPWR),
    .Y(_1650_),
    .VSS(VGND),
    .A1(net1088),
    .A2(net628));
 sg13g2_nand2_1 _4704_ (.Y(_1651_),
    .A(net731),
    .B(net715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4705_ (.Y(_1652_),
    .A(net711),
    .B(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4706_ (.Y(_1653_),
    .A(net738),
    .B(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or2_1 _4707_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1654_),
    .B(_1653_),
    .A(_1652_));
 sg13g2_o21ai_1 _4708_ (.B1(_1654_),
    .VDD(VPWR),
    .Y(_1655_),
    .VSS(VGND),
    .A1(net749),
    .A2(_1592_));
 sg13g2_xor2_1 _4709_ (.B(_1655_),
    .A(_1595_),
    .X(_1656_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4710_ (.Y(_1657_),
    .B(_1656_),
    .A_N(_1651_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4711_ (.B(_1656_),
    .A(_1651_),
    .X(_1658_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4712_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1591_),
    .A2(_1599_),
    .Y(_1659_),
    .B1(_1598_));
 sg13g2_nor2_1 _4713_ (.A(_1658_),
    .B(_1659_),
    .Y(_1660_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4714_ (.Y(_1661_),
    .A(_1658_),
    .B(_1659_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4715_ (.B(_1605_),
    .C(_1661_),
    .A(_1602_),
    .Y(_1662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4716_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1602_),
    .A2(_1605_),
    .Y(_1663_),
    .B1(_1661_));
 sg13g2_nand2_1 _4717_ (.Y(_1664_),
    .A(_1309_),
    .B(_1662_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4718_ (.A(net747),
    .B(net565),
    .Y(_1665_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4719_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2297_),
    .A2(net565),
    .Y(_1666_),
    .B1(_1665_));
 sg13g2_nor2_1 _4720_ (.A(_1246_),
    .B(_1273_),
    .Y(_1667_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4721_ (.Y(_1668_),
    .A(_1247_),
    .B(_1273_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4722_ (.B1(_1215_),
    .VDD(VPWR),
    .Y(_1669_),
    .VSS(VGND),
    .A1(_1218_),
    .A2(_1611_));
 sg13g2_xnor2_1 _4723_ (.Y(_1670_),
    .A(_1246_),
    .B(_1669_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4724_ (.B1(_1323_),
    .VDD(VPWR),
    .Y(_1671_),
    .VSS(VGND),
    .A1(net748),
    .A2(_1325_));
 sg13g2_a21oi_1 _4725_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1244_),
    .A2(_1383_),
    .Y(_1672_),
    .B1(_1313_));
 sg13g2_a21oi_1 _4726_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1243_),
    .A2(_1319_),
    .Y(_1673_),
    .B1(_1299_));
 sg13g2_o21ai_1 _4727_ (.B1(_1673_),
    .VDD(VPWR),
    .Y(_1674_),
    .VSS(VGND),
    .A1(_1245_),
    .A2(_1672_));
 sg13g2_a221oi_1 _4728_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1247_),
    .C1(_1674_),
    .B1(_1671_),
    .A1(_1244_),
    .Y(_1675_),
    .A2(_1327_));
 sg13g2_o21ai_1 _4729_ (.B1(_1675_),
    .VDD(VPWR),
    .Y(_1676_),
    .VSS(VGND),
    .A1(_1374_),
    .A2(_1670_));
 sg13g2_a221oi_1 _4730_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net631),
    .C1(_1676_),
    .B1(_1668_),
    .A1(net616),
    .Y(_1677_),
    .A2(_1666_));
 sg13g2_nand3b_1 _4731_ (.B(_1565_),
    .C(_1638_),
    .Y(_1678_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1494_));
 sg13g2_o21ai_1 _4732_ (.B1(_1678_),
    .VDD(VPWR),
    .Y(_1679_),
    .VSS(VGND),
    .A1(_1567_),
    .A2(_1640_));
 sg13g2_nand2b_1 _4733_ (.Y(_1680_),
    .B(_1638_),
    .A_N(_1563_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4734_ (.B1(_1636_),
    .VDD(VPWR),
    .Y(_1681_),
    .VSS(VGND),
    .A1(_1550_),
    .A2(_1637_));
 sg13g2_or2_1 _4735_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1682_),
    .B(_1625_),
    .A(_1623_));
 sg13g2_nand2_1 _4736_ (.Y(_1683_),
    .A(net746),
    .B(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4737_ (.Y(_1684_),
    .B(_1682_),
    .A_N(_1683_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4738_ (.B(_1683_),
    .A(_1682_),
    .X(_1685_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4739_ (.B1(_1633_),
    .VDD(VPWR),
    .Y(_1686_),
    .VSS(VGND),
    .A1(_1627_),
    .A2(_1634_));
 sg13g2_nand2_1 _4740_ (.Y(_1687_),
    .A(net742),
    .B(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4741_ (.A(net719),
    .B(net769),
    .X(_1688_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4742_ (.Y(_1689_),
    .B(_1688_),
    .A_N(_1529_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4743_ (.B(_1688_),
    .A(_1529_),
    .X(_1690_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4744_ (.B(_1690_),
    .A(_1687_),
    .X(_1691_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4745_ (.B1(_1629_),
    .VDD(VPWR),
    .Y(_1692_),
    .VSS(VGND),
    .A1(_1392_),
    .A2(_1630_));
 sg13g2_nand2_1 _4746_ (.Y(_1693_),
    .A(net723),
    .B(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4747_ (.A(net732),
    .B(net728),
    .C(net762),
    .D(net756),
    .X(_1694_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4748_ (.B(net728),
    .C(net762),
    .A(net732),
    .Y(_1695_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net756));
 sg13g2_a22oi_1 _4749_ (.Y(_1696_),
    .B1(net757),
    .B2(net733),
    .A2(net762),
    .A1(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _4750_ (.A(_1693_),
    .B(_1694_),
    .C(_1696_),
    .X(_1697_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4751_ (.B1(_1693_),
    .VDD(VPWR),
    .Y(_1698_),
    .VSS(VGND),
    .A1(_1694_),
    .A2(_1696_));
 sg13g2_nand3_1 _4752_ (.B(_1697_),
    .C(_1698_),
    .A(_1692_),
    .Y(_1699_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4753_ (.A2(_1698_),
    .A1(_1697_),
    .B1(_1692_),
    .X(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4754_ (.Y(_1701_),
    .A(_1699_),
    .B(_1700_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4755_ (.B(_1699_),
    .C(_1700_),
    .A(_1691_),
    .Y(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4756_ (.B(_1701_),
    .A(_1691_),
    .X(_1703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4757_ (.Y(_1704_),
    .B(_1686_),
    .A_N(_1703_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4758_ (.A(_1686_),
    .B_N(_1703_),
    .Y(_1705_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4759_ (.B(_1703_),
    .A(_1686_),
    .X(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4760_ (.Y(_1707_),
    .A(_1685_),
    .B(_1706_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4761_ (.Y(_1708_),
    .B(_1681_),
    .A_N(_1707_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4762_ (.B(_1707_),
    .A(_1681_),
    .X(_1709_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4763_ (.A(_1680_),
    .B(_1709_),
    .Y(_1710_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4764_ (.B(_1709_),
    .A(_1680_),
    .X(_1711_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4765_ (.B1(net615),
    .VDD(VPWR),
    .Y(_1712_),
    .VSS(VGND),
    .A1(_1679_),
    .A2(_1711_));
 sg13g2_a21o_2 _4766_ (.A2(_1711_),
    .A1(_1679_),
    .B1(_1712_),
    .X(_1713_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4767_ (.A(_1677_),
    .B(_1713_),
    .X(_1714_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4768_ (.B1(_1714_),
    .VDD(VPWR),
    .Y(_1715_),
    .VSS(VGND),
    .A1(_1663_),
    .A2(_1664_));
 sg13g2_nand2_1 _4769_ (.Y(_1716_),
    .A(_1404_),
    .B(_1646_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4770_ (.Y(_1717_),
    .A(net1037),
    .B(_1716_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4771_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net639),
    .C1(net630),
    .B1(_1717_),
    .A1(net614),
    .Y(_1718_),
    .A2(_1715_));
 sg13g2_nor2_1 _4772_ (.A(_1650_),
    .B(_1718_),
    .Y(_0301_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4773_ (.B1(_1657_),
    .VDD(VPWR),
    .Y(_1719_),
    .VSS(VGND),
    .A1(_1595_),
    .A2(_1655_));
 sg13g2_xnor2_1 _4774_ (.Y(_1720_),
    .A(net705),
    .B(_1654_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4775_ (.A(_1720_),
    .B_N(_1719_),
    .Y(_1721_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4776_ (.Y(_1722_),
    .A(_1719_),
    .B(_1720_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4777_ (.B1(_1722_),
    .VDD(VPWR),
    .Y(_1723_),
    .VSS(VGND),
    .A1(_1660_),
    .A2(_1663_));
 sg13g2_nor3_1 _4778_ (.A(_1660_),
    .B(_1663_),
    .C(_1722_),
    .Y(_1724_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4779_ (.A(_1310_),
    .B(_1724_),
    .Y(_1725_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4780_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1246_),
    .A2(_1669_),
    .Y(_1726_),
    .B1(_1243_));
 sg13g2_o21ai_1 _4781_ (.B1(_1373_),
    .VDD(VPWR),
    .Y(_1727_),
    .VSS(VGND),
    .A1(net632),
    .A2(_1726_));
 sg13g2_a21oi_1 _4782_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1242_),
    .A2(_1726_),
    .Y(_1728_),
    .B1(_1727_));
 sg13g2_nor2b_1 _4783_ (.A(net720),
    .B_N(net747),
    .Y(_1729_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4784_ (.A(net632),
    .B(_1667_),
    .C(_1729_),
    .Y(_1730_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4785_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net632),
    .A2(net565),
    .Y(_1731_),
    .B1(_1730_));
 sg13g2_nand2_1 _4786_ (.Y(_1732_),
    .A(net631),
    .B(_1731_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4787_ (.Y(_1733_),
    .A(_1240_),
    .B(_1324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4788_ (.B1(_1733_),
    .VDD(VPWR),
    .Y(_1734_),
    .VSS(VGND),
    .A1(_1240_),
    .A2(_1314_));
 sg13g2_nor2_1 _4789_ (.A(net632),
    .B(_1383_),
    .Y(_1735_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4790_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1242_),
    .A2(_1323_),
    .Y(_1736_),
    .B1(_1735_));
 sg13g2_mux2_1 _4791_ (.A0(_1280_),
    .A1(_1327_),
    .S(_1241_),
    .X(_1737_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor4_1 _4792_ (.A(_1728_),
    .B(_1734_),
    .C(_1736_),
    .D(_1737_),
    .Y(_1738_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4793_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1679_),
    .A2(_1711_),
    .Y(_1739_),
    .B1(_1710_));
 sg13g2_o21ai_1 _4794_ (.B1(_1704_),
    .VDD(VPWR),
    .Y(_1740_),
    .VSS(VGND),
    .A1(_1685_),
    .A2(_1705_));
 sg13g2_o21ai_1 _4795_ (.B1(_1689_),
    .VDD(VPWR),
    .Y(_1741_),
    .VSS(VGND),
    .A1(_1687_),
    .A2(_1690_));
 sg13g2_nor2_1 _4796_ (.A(net746),
    .B(net706),
    .Y(_1742_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4797_ (.A(_1653_),
    .B(_1687_),
    .Y(_1743_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4798_ (.Y(_1744_),
    .B1(net751),
    .B2(net738),
    .A2(net748),
    .A1(net742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4799_ (.A(_1743_),
    .B(_1744_),
    .Y(_1745_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4800_ (.B(_1745_),
    .A(_1742_),
    .X(_1746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4801_ (.Y(_1747_),
    .A(_1741_),
    .B(_1746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4802_ (.Y(_1748_),
    .A(_1741_),
    .B(_1746_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4803_ (.Y(_1749_),
    .A(_1699_),
    .B(_1702_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4804_ (.Y(_1750_),
    .A(net732),
    .B(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _4805_ (.A(net713),
    .B(net766),
    .X(_1751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _4806_ (.Y(_1752_),
    .A(net711),
    .B(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4807_ (.Y(_1753_),
    .A(net713),
    .B(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4808_ (.Y(_1754_),
    .A(_1688_),
    .B(_1751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4809_ (.Y(_1755_),
    .B1(net766),
    .B2(net719),
    .A2(net768),
    .A1(net713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4810_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1688_),
    .A2(_1751_),
    .Y(_1756_),
    .B1(_1755_));
 sg13g2_xor2_1 _4811_ (.B(_1756_),
    .A(_1750_),
    .X(_1757_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4812_ (.B1(_1695_),
    .VDD(VPWR),
    .Y(_1758_),
    .VSS(VGND),
    .A1(_1693_),
    .A2(_1696_));
 sg13g2_nand2_1 _4813_ (.Y(_1759_),
    .A(net723),
    .B(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4814_ (.X(_1760_),
    .A(net728),
    .B(\falu_i.falutop.alu_data_in[7] ),
    .C(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4815_ (.B(\falu_i.falutop.alu_data_in[7] ),
    .C(net755),
    .A(net727),
    .Y(_1761_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4816_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net728),
    .A2(net758),
    .Y(_1762_),
    .B1(\falu_i.falutop.alu_data_in[7] ));
 sg13g2_or3_1 _4817_ (.A(_1759_),
    .B(_1760_),
    .C(_1762_),
    .X(_1763_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4818_ (.B1(_1759_),
    .VDD(VPWR),
    .Y(_1764_),
    .VSS(VGND),
    .A1(_1760_),
    .A2(_1762_));
 sg13g2_nand3_1 _4819_ (.B(_1763_),
    .C(_1764_),
    .A(_1758_),
    .Y(_1765_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4820_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1763_),
    .A2(_1764_),
    .Y(_1766_),
    .B1(_1758_));
 sg13g2_a21o_1 _4821_ (.A2(_1764_),
    .A1(_1763_),
    .B1(_1758_),
    .X(_1767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4822_ (.Y(_1768_),
    .A(_1765_),
    .B(_1767_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4823_ (.Y(_1769_),
    .A(_1757_),
    .B(_1768_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4824_ (.Y(_1770_),
    .B(_1749_),
    .A_N(_1769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4825_ (.A(_1749_),
    .B_N(_1769_),
    .Y(_1771_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4826_ (.Y(_1772_),
    .A(_1749_),
    .B(_1769_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4827_ (.Y(_1773_),
    .A(_1748_),
    .B(_1772_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4828_ (.Y(_1774_),
    .A(_1740_),
    .B(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4829_ (.Y(_1775_),
    .A(_1740_),
    .B(_1773_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4830_ (.B(_1775_),
    .A(_1684_),
    .X(_1776_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4831_ (.Y(_1777_),
    .B(_1776_),
    .A_N(_1708_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4832_ (.B(_1776_),
    .A(_1708_),
    .X(_1778_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4833_ (.B(_1778_),
    .A(_1739_),
    .X(_1779_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4834_ (.Y(_1780_),
    .B1(_1779_),
    .B2(net615),
    .A2(_1725_),
    .A1(_1723_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4835_ (.B(_1738_),
    .C(_1780_),
    .A(_1732_),
    .Y(_1781_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4836_ (.B1(_1404_),
    .VDD(VPWR),
    .Y(_1782_),
    .VSS(VGND),
    .A1(net1037),
    .A2(_1646_));
 sg13g2_xnor2_1 _4837_ (.Y(_1783_),
    .A(\falu_i.falutop.div_inst.val[7] ),
    .B(_1782_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4838_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net639),
    .C1(_1075_),
    .B1(_1783_),
    .A1(net614),
    .Y(_1784_),
    .A2(_1781_));
 sg13g2_o21ai_1 _4839_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1785_),
    .VSS(VGND),
    .A1(net1041),
    .A2(net628));
 sg13g2_nor2_1 _4840_ (.A(_1784_),
    .B(_1785_),
    .Y(_0302_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4841_ (.B1(_1723_),
    .VDD(VPWR),
    .Y(_1786_),
    .VSS(VGND),
    .A1(net705),
    .A2(_1654_));
 sg13g2_o21ai_1 _4842_ (.B1(_1309_),
    .VDD(VPWR),
    .Y(_1787_),
    .VSS(VGND),
    .A1(_1721_),
    .A2(_1786_));
 sg13g2_o21ai_1 _4843_ (.B1(_1777_),
    .VDD(VPWR),
    .Y(_1788_),
    .VSS(VGND),
    .A1(_1739_),
    .A2(_1778_));
 sg13g2_o21ai_1 _4844_ (.B1(_1774_),
    .VDD(VPWR),
    .Y(_1789_),
    .VSS(VGND),
    .A1(_1684_),
    .A2(_1775_));
 sg13g2_o21ai_1 _4845_ (.B1(_1770_),
    .VDD(VPWR),
    .Y(_1790_),
    .VSS(VGND),
    .A1(_1748_),
    .A2(_1771_));
 sg13g2_a21oi_1 _4846_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1742_),
    .A2(_1745_),
    .Y(_1791_),
    .B1(_1743_));
 sg13g2_o21ai_1 _4847_ (.B1(_1754_),
    .VDD(VPWR),
    .Y(_1792_),
    .VSS(VGND),
    .A1(_1750_),
    .A2(_1755_));
 sg13g2_nor2_1 _4848_ (.A(net742),
    .B(net706),
    .Y(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4849_ (.A(net742),
    .B(net706),
    .C(_1653_),
    .Y(_1794_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _4850_ (.VDD(VPWR),
    .Y(_1795_),
    .A(_1794_),
    .VSS(VGND));
 sg13g2_xnor2_1 _4851_ (.Y(_1796_),
    .A(_1653_),
    .B(_1793_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4852_ (.Y(_1797_),
    .A(_1792_),
    .B(_1796_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4853_ (.A(_1791_),
    .B(_1797_),
    .Y(_1798_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4854_ (.Y(_1799_),
    .A(_1791_),
    .B(_1797_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4855_ (.B1(_1765_),
    .VDD(VPWR),
    .Y(_1800_),
    .VSS(VGND),
    .A1(_1757_),
    .A2(_1766_));
 sg13g2_nand2_1 _4856_ (.Y(_1801_),
    .A(net733),
    .B(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4857_ (.Y(_1802_),
    .B1(net752),
    .B2(net727),
    .A2(net768),
    .A1(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _4858_ (.X(_1803_),
    .A(net711),
    .B(net768),
    .C(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4859_ (.B(net768),
    .C(net752),
    .A(net711),
    .Y(_1804_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4860_ (.Y(_1805_),
    .A(net727),
    .B(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4861_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net727),
    .A2(_1803_),
    .Y(_1806_),
    .B1(_1802_));
 sg13g2_xor2_1 _4862_ (.B(_1806_),
    .A(_1801_),
    .X(_1807_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4863_ (.B1(_1761_),
    .VDD(VPWR),
    .Y(_1808_),
    .VSS(VGND),
    .A1(_1759_),
    .A2(_1762_));
 sg13g2_and4_1 _4864_ (.A(net723),
    .B(net718),
    .C(net761),
    .D(net755),
    .X(_1809_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _4865_ (.B(net718),
    .C(net761),
    .A(net723),
    .Y(_1810_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(net755));
 sg13g2_a22oi_1 _4866_ (.Y(_1811_),
    .B1(net755),
    .B2(net723),
    .A2(net761),
    .A1(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _4867_ (.B(_1751_),
    .C(_1810_),
    .Y(_1812_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1811_));
 sg13g2_o21ai_1 _4868_ (.B1(_1752_),
    .VDD(VPWR),
    .Y(_1813_),
    .VSS(VGND),
    .A1(_1809_),
    .A2(_1811_));
 sg13g2_and3_1 _4869_ (.X(_1814_),
    .A(_1808_),
    .B(_1812_),
    .C(_1813_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4870_ (.B(_1812_),
    .C(_1813_),
    .A(_1808_),
    .Y(_1815_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4871_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1812_),
    .A2(_1813_),
    .Y(_1816_),
    .B1(_1808_));
 sg13g2_or3_1 _4872_ (.A(_1807_),
    .B(_1814_),
    .C(_1816_),
    .X(_1817_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4873_ (.B1(_1807_),
    .VDD(VPWR),
    .Y(_1818_),
    .VSS(VGND),
    .A1(_1814_),
    .A2(_1816_));
 sg13g2_and3_1 _4874_ (.X(_1819_),
    .A(_1800_),
    .B(_1817_),
    .C(_1818_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4875_ (.B(_1817_),
    .C(_1818_),
    .A(_1800_),
    .Y(_1820_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4876_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1817_),
    .A2(_1818_),
    .Y(_1821_),
    .B1(_1800_));
 sg13g2_nor2_1 _4877_ (.A(_1819_),
    .B(_1821_),
    .Y(_1822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4878_ (.Y(_1823_),
    .A(_1799_),
    .B(_1822_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4879_ (.Y(_1824_),
    .A(_1790_),
    .B(_1823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4880_ (.Y(_1825_),
    .A(_1790_),
    .B(_1823_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4881_ (.B(_1825_),
    .A(_1747_),
    .X(_1826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4882_ (.Y(_1827_),
    .A(_1789_),
    .B(_1826_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4883_ (.B(_1826_),
    .A(_1789_),
    .X(_1828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4884_ (.Y(_1829_),
    .A(_1788_),
    .B(_1828_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4885_ (.B1(net615),
    .VDD(VPWR),
    .Y(_1830_),
    .VSS(VGND),
    .A1(_1788_),
    .A2(_1828_));
 sg13g2_nand2b_2 _4886_ (.Y(_1831_),
    .B(_1829_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1830_));
 sg13g2_nor2_1 _4887_ (.A(_1240_),
    .B(_1727_),
    .Y(_1832_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4888_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net632),
    .A2(net565),
    .Y(_1833_),
    .B1(_1276_));
 sg13g2_a21oi_2 _4889_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1832_),
    .Y(_1834_),
    .A2(_1833_),
    .A1(net631));
 sg13g2_a21oi_1 _4890_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2301_),
    .A2(net564),
    .Y(_1835_),
    .B1(_1282_));
 sg13g2_o21ai_1 _4891_ (.B1(_1835_),
    .VDD(VPWR),
    .Y(_1836_),
    .VSS(VGND),
    .A1(net744),
    .A2(net563));
 sg13g2_nand4_1 _4892_ (.B(_1831_),
    .C(_1834_),
    .A(_1787_),
    .Y(_1837_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_1836_));
 sg13g2_a221oi_1 _4893_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1837_),
    .C1(net630),
    .B1(net614),
    .A1(\falu_i.falutop.div_inst.rem[0] ),
    .Y(_1838_),
    .A2(net638));
 sg13g2_o21ai_1 _4894_ (.B1(net815),
    .VDD(VPWR),
    .Y(_1839_),
    .VSS(VGND),
    .A1(net1033),
    .A2(net627));
 sg13g2_nor2_1 _4895_ (.A(_1838_),
    .B(_1839_),
    .Y(_0303_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4896_ (.B1(net815),
    .VDD(VPWR),
    .Y(_1840_),
    .VSS(VGND),
    .A1(net1064),
    .A2(net627));
 sg13g2_o21ai_1 _4897_ (.B1(_1824_),
    .VDD(VPWR),
    .Y(_1841_),
    .VSS(VGND),
    .A1(_1747_),
    .A2(_1825_));
 sg13g2_a21oi_1 _4898_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1792_),
    .A2(_1796_),
    .Y(_1842_),
    .B1(_1798_));
 sg13g2_o21ai_1 _4899_ (.B1(_1820_),
    .VDD(VPWR),
    .Y(_1843_),
    .VSS(VGND),
    .A1(_1799_),
    .A2(_1821_));
 sg13g2_o21ai_1 _4900_ (.B1(_1805_),
    .VDD(VPWR),
    .Y(_1844_),
    .VSS(VGND),
    .A1(_1801_),
    .A2(_1802_));
 sg13g2_nand2_1 _4901_ (.Y(_1845_),
    .A(net733),
    .B(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4902_ (.A(net738),
    .B(net706),
    .Y(_1846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4903_ (.Y(_1847_),
    .B(_1846_),
    .A_N(_1845_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4904_ (.Y(_1848_),
    .A(_1845_),
    .B(_1846_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4905_ (.Y(_1849_),
    .A(_1844_),
    .B(_1848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4906_ (.Y(_1850_),
    .A(_1844_),
    .B(_1848_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4907_ (.Y(_1851_),
    .A(_1795_),
    .B(_1850_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4908_ (.B1(_1815_),
    .VDD(VPWR),
    .Y(_1852_),
    .VSS(VGND),
    .A1(_1807_),
    .A2(_1816_));
 sg13g2_nand2_1 _4909_ (.Y(_1853_),
    .A(net727),
    .B(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4910_ (.Y(_1854_),
    .A(net723),
    .B(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4911_ (.Y(_1855_),
    .A(_1622_),
    .B(_1753_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4912_ (.Y(_1856_),
    .A(_1853_),
    .B(_1855_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4913_ (.B1(_1810_),
    .VDD(VPWR),
    .Y(_1857_),
    .VSS(VGND),
    .A1(_1752_),
    .A2(_1811_));
 sg13g2_a22oi_1 _4914_ (.Y(_1858_),
    .B1(net758),
    .B2(net718),
    .A2(net761),
    .A1(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _4915_ (.A(net719),
    .B(net712),
    .C(net761),
    .D(net758),
    .X(_1859_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4916_ (.B1(_1752_),
    .VDD(VPWR),
    .Y(_1860_),
    .VSS(VGND),
    .A1(_1858_),
    .A2(_1859_));
 sg13g2_or3_1 _4917_ (.A(_1752_),
    .B(_1858_),
    .C(_1859_),
    .X(_1861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_1 _4918_ (.X(_1862_),
    .A(_1857_),
    .B(_1860_),
    .C(_1861_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4919_ (.B(_1860_),
    .C(_1861_),
    .A(_1857_),
    .Y(_1863_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4920_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1860_),
    .A2(_1861_),
    .Y(_1864_),
    .B1(_1857_));
 sg13g2_or3_1 _4921_ (.A(_1856_),
    .B(_1862_),
    .C(_1864_),
    .X(_1865_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4922_ (.B1(_1856_),
    .VDD(VPWR),
    .Y(_1866_),
    .VSS(VGND),
    .A1(_1862_),
    .A2(_1864_));
 sg13g2_and3_1 _4923_ (.X(_1867_),
    .A(_1852_),
    .B(_1865_),
    .C(_1866_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4924_ (.B(_1865_),
    .C(_1866_),
    .A(_1852_),
    .Y(_1868_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4925_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1865_),
    .A2(_1866_),
    .Y(_1869_),
    .B1(_1852_));
 sg13g2_or3_1 _4926_ (.A(_1851_),
    .B(_1867_),
    .C(_1869_),
    .X(_1870_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4927_ (.B1(_1851_),
    .VDD(VPWR),
    .Y(_1871_),
    .VSS(VGND),
    .A1(_1867_),
    .A2(_1869_));
 sg13g2_nand3_1 _4928_ (.B(_1870_),
    .C(_1871_),
    .A(_1843_),
    .Y(_1872_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4929_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1870_),
    .A2(_1871_),
    .Y(_1873_),
    .B1(_1843_));
 sg13g2_a21o_1 _4930_ (.A2(_1871_),
    .A1(_1870_),
    .B1(_1843_),
    .X(_1874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4931_ (.Y(_1875_),
    .A(_1872_),
    .B(_1874_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4932_ (.Y(_1876_),
    .A(_1842_),
    .B(_1875_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4933_ (.A(_1841_),
    .B_N(_1876_),
    .Y(_1877_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4934_ (.Y(_1878_),
    .B(_1841_),
    .A_N(_1876_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4935_ (.B(_1876_),
    .A(_1841_),
    .X(_1879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _4936_ (.A2(_1829_),
    .A1(_1827_),
    .B1(_1879_),
    .X(_1880_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4937_ (.B(_1829_),
    .C(_1879_),
    .A(_1827_),
    .Y(_1881_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4938_ (.B(_1880_),
    .C(_1881_),
    .A(_1317_),
    .Y(_1882_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4939_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2304_),
    .A2(net563),
    .Y(_1883_),
    .B1(_1282_));
 sg13g2_o21ai_1 _4940_ (.B1(_1883_),
    .VDD(VPWR),
    .Y(_1884_),
    .VSS(VGND),
    .A1(net740),
    .A2(net564));
 sg13g2_nand3_1 _4941_ (.B(_1882_),
    .C(_1884_),
    .A(_1834_),
    .Y(_1885_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _4942_ (.B(\falu_i.falutop.div_inst.rem[1] ),
    .C(\falu_i.falutop.div_inst.rem[0] ),
    .A(net775),
    .Y(_1886_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4943_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net775),
    .A2(\falu_i.falutop.div_inst.rem[0] ),
    .Y(_1887_),
    .B1(\falu_i.falutop.div_inst.rem[1] ));
 sg13g2_nor2_1 _4944_ (.A(_1074_),
    .B(_1887_),
    .Y(_1888_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4945_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1888_),
    .C1(net630),
    .B1(_1886_),
    .A1(net614),
    .Y(_1889_),
    .A2(_1885_));
 sg13g2_nor2_1 _4946_ (.A(_1840_),
    .B(_1889_),
    .Y(_0304_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4947_ (.B1(_1872_),
    .VDD(VPWR),
    .Y(_1890_),
    .VSS(VGND),
    .A1(_1842_),
    .A2(_1873_));
 sg13g2_o21ai_1 _4948_ (.B1(_1849_),
    .VDD(VPWR),
    .Y(_1891_),
    .VSS(VGND),
    .A1(_1795_),
    .A2(_1850_));
 sg13g2_inv_1 _4949_ (.VDD(VPWR),
    .Y(_1892_),
    .A(_1891_),
    .VSS(VGND));
 sg13g2_o21ai_1 _4950_ (.B1(_1868_),
    .VDD(VPWR),
    .Y(_1893_),
    .VSS(VGND),
    .A1(_1851_),
    .A2(_1869_));
 sg13g2_o21ai_1 _4951_ (.B1(_1854_),
    .VDD(VPWR),
    .Y(_1894_),
    .VSS(VGND),
    .A1(_1853_),
    .A2(_1855_));
 sg13g2_nand2_1 _4952_ (.Y(_1895_),
    .A(net727),
    .B(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4953_ (.A(net733),
    .B(net705),
    .Y(_1896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4954_ (.Y(_1897_),
    .B(_1896_),
    .A_N(_1895_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4955_ (.Y(_1898_),
    .A(_1895_),
    .B(_1896_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4956_ (.Y(_1899_),
    .A(_1894_),
    .B(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4957_ (.Y(_1900_),
    .A(_1894_),
    .B(_1898_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4958_ (.Y(_1901_),
    .A(_1847_),
    .B(_1900_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4959_ (.B1(_1863_),
    .VDD(VPWR),
    .Y(_1902_),
    .VSS(VGND),
    .A1(_1856_),
    .A2(_1864_));
 sg13g2_nand2_1 _4960_ (.Y(_1903_),
    .A(net718),
    .B(_1803_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4961_ (.Y(_1904_),
    .B1(net753),
    .B2(net718),
    .A2(net768),
    .A1(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4962_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net718),
    .A2(_1803_),
    .Y(_1905_),
    .B1(_1904_));
 sg13g2_xnor2_1 _4963_ (.Y(_1906_),
    .A(_1214_),
    .B(_1905_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4964_ (.B1(net712),
    .VDD(VPWR),
    .Y(_1907_),
    .VSS(VGND),
    .A1(net761),
    .A2(net755));
 sg13g2_nand3_1 _4965_ (.B(net764),
    .C(net755),
    .A(net711),
    .Y(_1908_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _4966_ (.Y(_1909_),
    .B(_1908_),
    .A_N(_1907_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _4967_ (.Y(_1910_),
    .B1(_1859_),
    .B2(_2304_),
    .A2(_1858_),
    .A1(_1751_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4968_ (.Y(_1911_),
    .A(_1909_),
    .B(_1910_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4969_ (.B(_1911_),
    .A(_1906_),
    .X(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4970_ (.Y(_1913_),
    .A(_1902_),
    .B(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4971_ (.Y(_1914_),
    .A(_1902_),
    .B(_1912_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4972_ (.B(_1914_),
    .A(_1901_),
    .X(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4973_ (.Y(_1916_),
    .A(_1893_),
    .B(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4974_ (.Y(_1917_),
    .A(_1893_),
    .B(_1915_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4975_ (.Y(_1918_),
    .A(_1892_),
    .B(_1917_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4976_ (.A(_1918_),
    .B_N(_1890_),
    .Y(_1919_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _4977_ (.B(_1918_),
    .A(_1890_),
    .X(_1920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _4978_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1878_),
    .A2(_1880_),
    .Y(_1921_),
    .B1(_1920_));
 sg13g2_and3_1 _4979_ (.X(_1922_),
    .A(_1878_),
    .B(_1880_),
    .C(_1920_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_2 _4980_ (.A(_1318_),
    .B(_1921_),
    .C(_1922_),
    .Y(_1923_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _4981_ (.A(net765),
    .B_N(net563),
    .Y(_1924_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4982_ (.B1(net616),
    .VDD(VPWR),
    .Y(_1925_),
    .VSS(VGND),
    .A1(net739),
    .A2(net563));
 sg13g2_o21ai_1 _4983_ (.B1(_1834_),
    .VDD(VPWR),
    .Y(_1926_),
    .VSS(VGND),
    .A1(_1924_),
    .A2(_1925_));
 sg13g2_or2_1 _4984_ (.VSS(VGND),
    .VDD(VPWR),
    .X(_1927_),
    .B(_1926_),
    .A(_1923_));
 sg13g2_o21ai_1 _4985_ (.B1(net774),
    .VDD(VPWR),
    .Y(_1928_),
    .VSS(VGND),
    .A1(\falu_i.falutop.div_inst.rem[1] ),
    .A2(\falu_i.falutop.div_inst.rem[0] ));
 sg13g2_nand2b_1 _4986_ (.Y(_1929_),
    .B(_1928_),
    .A_N(\falu_i.falutop.div_inst.rem[2] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4987_ (.Y(_1930_),
    .A(\falu_i.falutop.div_inst.rem[2] ),
    .B(_1928_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _4988_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net638),
    .C1(net630),
    .B1(_1930_),
    .A1(net614),
    .Y(_1931_),
    .A2(_1927_));
 sg13g2_o21ai_1 _4989_ (.B1(net818),
    .VDD(VPWR),
    .Y(_1932_),
    .VSS(VGND),
    .A1(net1062),
    .A2(net629));
 sg13g2_nor2_1 _4990_ (.A(_1931_),
    .B(_1932_),
    .Y(_0305_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _4991_ (.B1(_1916_),
    .VDD(VPWR),
    .Y(_1933_),
    .VSS(VGND),
    .A1(_1892_),
    .A2(_1917_));
 sg13g2_o21ai_1 _4992_ (.B1(_1899_),
    .VDD(VPWR),
    .Y(_1934_),
    .VSS(VGND),
    .A1(_1847_),
    .A2(_1900_));
 sg13g2_o21ai_1 _4993_ (.B1(_1913_),
    .VDD(VPWR),
    .Y(_1935_),
    .VSS(VGND),
    .A1(_1901_),
    .A2(_1914_));
 sg13g2_o21ai_1 _4994_ (.B1(_1903_),
    .VDD(VPWR),
    .Y(_1936_),
    .VSS(VGND),
    .A1(_1215_),
    .A2(_1904_));
 sg13g2_nand2_1 _4995_ (.Y(_1937_),
    .A(net723),
    .B(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _4996_ (.A(net727),
    .B(net705),
    .Y(_1938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _4997_ (.A(net727),
    .B(net706),
    .C(_1937_),
    .Y(_1939_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _4998_ (.Y(_1940_),
    .A(_1937_),
    .B(_1938_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _4999_ (.Y(_1941_),
    .A(_1936_),
    .B(_1940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5000_ (.Y(_1942_),
    .A(_1936_),
    .B(_1940_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5001_ (.Y(_1943_),
    .A(_1897_),
    .B(_1942_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and4_1 _5002_ (.A(net711),
    .B(net766),
    .C(net761),
    .D(net755),
    .X(_1944_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5003_ (.VDD(VPWR),
    .Y(_1945_),
    .A(_1944_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5004_ (.B1(_1945_),
    .VDD(VPWR),
    .Y(_1946_),
    .VSS(VGND),
    .A1(_1906_),
    .A2(_1911_));
 sg13g2_a21oi_2 _5005_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_1944_),
    .Y(_1947_),
    .A2(_1907_),
    .A1(_1752_));
 sg13g2_inv_1 _5006_ (.VDD(VPWR),
    .Y(_1948_),
    .A(_1947_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5007_ (.B1(net711),
    .VDD(VPWR),
    .Y(_1949_),
    .VSS(VGND),
    .A1(net768),
    .A2(net752));
 sg13g2_nor2_1 _5008_ (.A(_1803_),
    .B(_1949_),
    .Y(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5009_ (.Y(_1951_),
    .A(net718),
    .B(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5010_ (.A(_1803_),
    .B(_1949_),
    .C(_1951_),
    .Y(_1952_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5011_ (.B(_1951_),
    .A(_1950_),
    .X(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5012_ (.A(_1948_),
    .B(_1953_),
    .Y(_1954_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5013_ (.Y(_1955_),
    .A(_1948_),
    .B(_1953_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5014_ (.A(_1955_),
    .B_N(_1946_),
    .Y(_1956_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5015_ (.B(_1955_),
    .A(_1946_),
    .X(_1957_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5016_ (.A(_1943_),
    .B(_1957_),
    .Y(_1958_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5017_ (.B(_1957_),
    .A(_1943_),
    .X(_1959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5018_ (.Y(_1960_),
    .A(_1935_),
    .B(_1959_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5019_ (.A(_1960_),
    .B_N(_1934_),
    .Y(_1961_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5020_ (.Y(_1962_),
    .A(_1934_),
    .B(_1960_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5021_ (.A(_1933_),
    .B(_1962_),
    .Y(_1963_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5022_ (.Y(_1964_),
    .A(_1933_),
    .B(_1962_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5023_ (.VDD(VPWR),
    .Y(_1965_),
    .A(_1964_),
    .VSS(VGND));
 sg13g2_o21ai_1 _5024_ (.B1(_1965_),
    .VDD(VPWR),
    .Y(_1966_),
    .VSS(VGND),
    .A1(_1919_),
    .A2(_1921_));
 sg13g2_or3_1 _5025_ (.A(_1919_),
    .B(_1921_),
    .C(_1965_),
    .X(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and3_2 _5026_ (.X(_1968_),
    .A(net615),
    .B(_1966_),
    .C(_1967_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5027_ (.Y(_1969_),
    .B(net563),
    .A_N(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5028_ (.B1(_1969_),
    .VDD(VPWR),
    .Y(_1970_),
    .VSS(VGND),
    .A1(net731),
    .A2(net563));
 sg13g2_o21ai_1 _5029_ (.B1(_1834_),
    .VDD(VPWR),
    .Y(_1971_),
    .VSS(VGND),
    .A1(_1282_),
    .A2(_1970_));
 sg13g2_o21ai_1 _5030_ (.B1(_1590_),
    .VDD(VPWR),
    .Y(_1972_),
    .VSS(VGND),
    .A1(_1968_),
    .A2(_1971_));
 sg13g2_a21o_1 _5031_ (.A2(_1929_),
    .A1(net773),
    .B1(\falu_i.falutop.div_inst.rem[3] ),
    .X(_1973_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5032_ (.B(\falu_i.falutop.div_inst.rem[3] ),
    .C(_1929_),
    .A(net773),
    .Y(_1974_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5033_ (.B(_1973_),
    .C(_1974_),
    .A(net638),
    .Y(_1975_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5034_ (.A(net627),
    .B(_1975_),
    .X(_1976_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5035_ (.B1(net815),
    .VDD(VPWR),
    .Y(_1977_),
    .VSS(VGND),
    .A1(net1020),
    .A2(net627));
 sg13g2_a21oi_1 _5036_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1972_),
    .A2(_1976_),
    .Y(_0306_),
    .B1(_1977_));
 sg13g2_nor2_1 _5037_ (.A(_1920_),
    .B(_1964_),
    .Y(_1978_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5038_ (.Y(_1979_),
    .B(_1978_),
    .A_N(_1879_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3b_1 _5039_ (.B(_1788_),
    .C(_1828_),
    .Y(_1980_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_1979_));
 sg13g2_o21ai_1 _5040_ (.B1(_1878_),
    .VDD(VPWR),
    .Y(_1981_),
    .VSS(VGND),
    .A1(_1827_),
    .A2(_1877_));
 sg13g2_nor2b_1 _5041_ (.A(_1963_),
    .B_N(_1919_),
    .Y(_1982_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5042_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(_1981_),
    .C1(_1982_),
    .B1(_1978_),
    .A1(_1933_),
    .Y(_1983_),
    .A2(_1962_));
 sg13g2_a21o_1 _5043_ (.A2(_1959_),
    .A1(_1935_),
    .B1(_1961_),
    .X(_1984_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5044_ (.B1(_1941_),
    .VDD(VPWR),
    .Y(_1985_),
    .VSS(VGND),
    .A1(_1897_),
    .A2(_1942_));
 sg13g2_nor2_1 _5045_ (.A(_1956_),
    .B(_1958_),
    .Y(_1986_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5046_ (.Y(_1987_),
    .A(_1652_),
    .B(_1950_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5047_ (.Y(_1988_),
    .A(_1947_),
    .B(_1987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5048_ (.A(_1944_),
    .B(_1954_),
    .Y(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5049_ (.A(_1988_),
    .B(_1989_),
    .Y(_1990_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5050_ (.Y(_1991_),
    .A(_1988_),
    .B(_1989_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5051_ (.A(_1803_),
    .B(_1952_),
    .Y(_1992_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5052_ (.A(net724),
    .B(net705),
    .Y(_1993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5053_ (.A(net724),
    .B(net705),
    .C(_1244_),
    .Y(_1994_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5054_ (.Y(_1995_),
    .A(_1244_),
    .B(_1993_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5055_ (.A(_1992_),
    .B_N(_1995_),
    .Y(_1996_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5056_ (.Y(_1997_),
    .A(_1992_),
    .B(_1995_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5057_ (.Y(_1998_),
    .A(_1939_),
    .B(_1997_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5058_ (.A(_1991_),
    .B(_1998_),
    .Y(_1999_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5059_ (.Y(_2000_),
    .A(_1991_),
    .B(_1998_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5060_ (.A(_1986_),
    .B(_2000_),
    .Y(_2001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5061_ (.Y(_2002_),
    .A(_1986_),
    .B(_2000_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5062_ (.Y(_2003_),
    .B(_2002_),
    .A_N(_2001_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5063_ (.B(_2003_),
    .A(_1985_),
    .X(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5064_ (.A(_2004_),
    .B_N(_1984_),
    .Y(_2005_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5065_ (.Y(_2006_),
    .A(_1984_),
    .B(_2004_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5066_ (.VDD(VPWR),
    .Y(_2007_),
    .A(_2006_),
    .VSS(VGND));
 sg13g2_nand3_1 _5067_ (.B(_1983_),
    .C(_2007_),
    .A(_1980_),
    .Y(_2008_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_2 _5068_ (.VSS(VGND),
    .VDD(VPWR),
    .B1(_2007_),
    .Y(_2009_),
    .A2(_1983_),
    .A1(_1980_));
 sg13g2_nand3b_1 _5069_ (.B(_1317_),
    .C(_2008_),
    .Y(_2010_),
    .VDD(VPWR),
    .VSS(VGND),
    .A_N(_2009_));
 sg13g2_a21oi_1 _5070_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2303_),
    .A2(net566),
    .Y(_2011_),
    .B1(_1282_));
 sg13g2_o21ai_1 _5071_ (.B1(_2011_),
    .VDD(VPWR),
    .Y(_2012_),
    .VSS(VGND),
    .A1(net726),
    .A2(net566));
 sg13g2_nand3_1 _5072_ (.B(_2010_),
    .C(_2012_),
    .A(_1834_),
    .Y(_2013_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5073_ (.A2(_1973_),
    .A1(net773),
    .B1(\falu_i.falutop.div_inst.rem[4] ),
    .X(_2014_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5074_ (.B(\falu_i.falutop.div_inst.rem[4] ),
    .C(_1973_),
    .A(net773),
    .Y(_2015_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5075_ (.A(_2014_),
    .B(_2015_),
    .X(_2016_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5076_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net638),
    .C1(net630),
    .B1(_2016_),
    .A1(net614),
    .Y(_2017_),
    .A2(_2013_));
 sg13g2_o21ai_1 _5077_ (.B1(net815),
    .VDD(VPWR),
    .Y(_2018_),
    .VSS(VGND),
    .A1(net1018),
    .A2(net627));
 sg13g2_nor2_1 _5078_ (.A(_2017_),
    .B(_2018_),
    .Y(_0307_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5079_ (.A2(_1997_),
    .A1(_1939_),
    .B1(_1996_),
    .X(_2019_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5080_ (.A(_1990_),
    .B(_1999_),
    .Y(_2020_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5081_ (.Y(_2021_),
    .A(_1944_),
    .B(_1987_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5082_ (.A(_1944_),
    .B(_1947_),
    .C(_1987_),
    .X(_2022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_2 _5083_ (.Y(_2023_),
    .A(_2021_),
    .B(_2022_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5084_ (.B1(_1804_),
    .VDD(VPWR),
    .Y(_2024_),
    .VSS(VGND),
    .A1(_1652_),
    .A2(_1949_));
 sg13g2_inv_1 _5085_ (.VDD(VPWR),
    .Y(_2025_),
    .A(_2024_),
    .VSS(VGND));
 sg13g2_nor2b_2 _5086_ (.A(_1241_),
    .B_N(_1729_),
    .Y(_2026_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5087_ (.VDD(VPWR),
    .Y(_2027_),
    .A(_2026_),
    .VSS(VGND));
 sg13g2_a22oi_1 _5088_ (.Y(_2028_),
    .B1(net747),
    .B2(net714),
    .A2(\falu_i.falutop.alu_data_in[7] ),
    .A1(_2297_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5089_ (.A(_2026_),
    .B(_2028_),
    .Y(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5090_ (.A(_2024_),
    .B(_2029_),
    .X(_2030_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5091_ (.Y(_2031_),
    .A(_2025_),
    .B(_2029_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5092_ (.Y(_2032_),
    .A(_1994_),
    .B(_2031_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5093_ (.Y(_2033_),
    .A(_2023_),
    .B(_2032_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5094_ (.A(_2020_),
    .B(_2033_),
    .Y(_2034_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5095_ (.Y(_2035_),
    .A(_2020_),
    .B(_2033_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5096_ (.B(_2033_),
    .A(_2020_),
    .X(_2036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5097_ (.Y(_2037_),
    .A(_2019_),
    .B(_2036_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5098_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1985_),
    .A2(_2002_),
    .Y(_2038_),
    .B1(_2001_));
 sg13g2_xor2_1 _5099_ (.B(_2038_),
    .A(_2037_),
    .X(_2039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_or3_1 _5100_ (.A(_2005_),
    .B(_2009_),
    .C(_2039_),
    .X(_2040_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5101_ (.Y(_2041_),
    .A(_2009_),
    .B(_2039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5102_ (.Y(_2042_),
    .A(_2005_),
    .B(_2039_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand4_1 _5103_ (.B(_2040_),
    .C(_2041_),
    .A(_1317_),
    .Y(_2043_),
    .VDD(VPWR),
    .VSS(VGND),
    .D(_2042_));
 sg13g2_a21oi_1 _5104_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2305_),
    .A2(net564),
    .Y(_2044_),
    .B1(_1282_));
 sg13g2_o21ai_1 _5105_ (.B1(_2044_),
    .VDD(VPWR),
    .Y(_2045_),
    .VSS(VGND),
    .A1(net722),
    .A2(net564));
 sg13g2_nand3_1 _5106_ (.B(_2043_),
    .C(_2045_),
    .A(_1834_),
    .Y(_2046_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21o_1 _5107_ (.A2(_2014_),
    .A1(net773),
    .B1(\falu_i.falutop.div_inst.rem[5] ),
    .X(_2047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand3_1 _5108_ (.B(\falu_i.falutop.div_inst.rem[5] ),
    .C(_2014_),
    .A(net773),
    .Y(_2048_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_and2_1 _5109_ (.A(_2047_),
    .B(_2048_),
    .X(_2049_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a221oi_1 _5110_ (.VDD(VPWR),
    .VSS(VGND),
    .B2(net638),
    .C1(net630),
    .B1(_2049_),
    .A1(net614),
    .Y(_2050_),
    .A2(_2046_));
 sg13g2_o21ai_1 _5111_ (.B1(net815),
    .VDD(VPWR),
    .Y(_2051_),
    .VSS(VGND),
    .A1(net1035),
    .A2(net627));
 sg13g2_nor2_1 _5112_ (.A(_2050_),
    .B(_2051_),
    .Y(_0308_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5113_ (.B1(_2042_),
    .VDD(VPWR),
    .Y(_2052_),
    .VSS(VGND),
    .A1(_2037_),
    .A2(_2038_));
 sg13g2_a21oi_1 _5114_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2009_),
    .A2(_2039_),
    .Y(_2053_),
    .B1(_2052_));
 sg13g2_a21oi_1 _5115_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_1994_),
    .A2(_2031_),
    .Y(_2054_),
    .B1(_2030_));
 sg13g2_o21ai_1 _5116_ (.B1(_2021_),
    .VDD(VPWR),
    .Y(_2055_),
    .VSS(VGND),
    .A1(_2023_),
    .A2(_2032_));
 sg13g2_a21oi_1 _5117_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net714),
    .A2(net747),
    .Y(_2056_),
    .B1(_1275_));
 sg13g2_xnor2_1 _5118_ (.Y(_2057_),
    .A(_2024_),
    .B(_2056_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5119_ (.A(_2026_),
    .B(_2057_),
    .Y(_2058_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5120_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2025_),
    .A2(_2026_),
    .Y(_2059_),
    .B1(_2058_));
 sg13g2_xnor2_1 _5121_ (.Y(_2060_),
    .A(_2023_),
    .B(_2059_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5122_ (.B(_2060_),
    .A(_2055_),
    .X(_2061_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5123_ (.A(_2054_),
    .B_N(_2061_),
    .Y(_2062_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5124_ (.B(_2061_),
    .A(_2054_),
    .X(_2063_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5125_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2019_),
    .A2(_2035_),
    .Y(_2064_),
    .B1(_2034_));
 sg13g2_xnor2_1 _5126_ (.Y(_2065_),
    .A(_2063_),
    .B(_2064_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5127_ (.B1(net615),
    .VDD(VPWR),
    .Y(_2066_),
    .VSS(VGND),
    .A1(_2053_),
    .A2(_2065_));
 sg13g2_a21oi_1 _5128_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2053_),
    .A2(_2065_),
    .Y(_2067_),
    .B1(_2066_));
 sg13g2_nor2b_1 _5129_ (.A(net749),
    .B_N(net563),
    .Y(_2068_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5130_ (.B1(_1281_),
    .VDD(VPWR),
    .Y(_2069_),
    .VSS(VGND),
    .A1(net717),
    .A2(net563));
 sg13g2_o21ai_1 _5131_ (.B1(_1834_),
    .VDD(VPWR),
    .Y(_2070_),
    .VSS(VGND),
    .A1(_2068_),
    .A2(_2069_));
 sg13g2_o21ai_1 _5132_ (.B1(_1590_),
    .VDD(VPWR),
    .Y(_2071_),
    .VSS(VGND),
    .A1(_2067_),
    .A2(_2070_));
 sg13g2_nand2_1 _5133_ (.Y(_2072_),
    .A(net773),
    .B(_2047_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5134_ (.Y(_2073_),
    .A(\falu_i.falutop.div_inst.rem[6] ),
    .B(_2072_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5135_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net638),
    .A2(_2073_),
    .Y(_2074_),
    .B1(net630));
 sg13g2_o21ai_1 _5136_ (.B1(net815),
    .VDD(VPWR),
    .Y(_2075_),
    .VSS(VGND),
    .A1(net1071),
    .A2(net627));
 sg13g2_a21oi_1 _5137_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2071_),
    .A2(_2074_),
    .Y(_0309_),
    .B1(_2075_));
 sg13g2_a21oi_1 _5138_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2055_),
    .A2(_2060_),
    .Y(_2076_),
    .B1(_2062_));
 sg13g2_o21ai_1 _5139_ (.B1(_2027_),
    .VDD(VPWR),
    .Y(_2077_),
    .VSS(VGND),
    .A1(_2025_),
    .A2(_2056_));
 sg13g2_mux2_1 _5140_ (.A0(_2022_),
    .A1(_2021_),
    .S(_2057_),
    .X(_2078_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5141_ (.B1(_2078_),
    .VDD(VPWR),
    .Y(_2079_),
    .VSS(VGND),
    .A1(_2023_),
    .A2(_2027_));
 sg13g2_mux2_1 _5142_ (.A0(_2078_),
    .A1(_2079_),
    .S(_2077_),
    .X(_2080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5143_ (.Y(_2081_),
    .A(_2076_),
    .B(_2080_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5144_ (.B1(_2081_),
    .VDD(VPWR),
    .Y(_2082_),
    .VSS(VGND),
    .A1(_2063_),
    .A2(_2064_));
 sg13g2_nor2_1 _5145_ (.A(_2066_),
    .B(_2082_),
    .Y(_2083_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5146_ (.B1(_1834_),
    .VDD(VPWR),
    .Y(_2084_),
    .VSS(VGND),
    .A1(_1240_),
    .A2(_1282_));
 sg13g2_o21ai_1 _5147_ (.B1(_1590_),
    .VDD(VPWR),
    .Y(_2085_),
    .VSS(VGND),
    .A1(_2083_),
    .A2(_2084_));
 sg13g2_o21ai_1 _5148_ (.B1(net774),
    .VDD(VPWR),
    .Y(_2086_),
    .VSS(VGND),
    .A1(\falu_i.falutop.div_inst.rem[6] ),
    .A2(_2047_));
 sg13g2_xnor2_1 _5149_ (.Y(_2087_),
    .A(\falu_i.falutop.div_inst.rem[7] ),
    .B(_2086_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5150_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net638),
    .A2(_2087_),
    .Y(_2088_),
    .B1(net630));
 sg13g2_o21ai_1 _5151_ (.B1(net815),
    .VDD(VPWR),
    .Y(_2089_),
    .VSS(VGND),
    .A1(net1029),
    .A2(net627));
 sg13g2_a21oi_1 _5152_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2085_),
    .A2(_2088_),
    .Y(_0310_),
    .B1(_2089_));
 sg13g2_nor3_1 _5153_ (.A(\falu_i.falutop.data_in[8] ),
    .B(\falu_i.falutop.data_in[9] ),
    .C(\falu_i.falutop.data_in[10] ),
    .Y(_2090_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5154_ (.A(\falu_i.falutop.data_in[11] ),
    .B_N(_2090_),
    .Y(_2091_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5155_ (.A(\falu_i.falutop.data_in[12] ),
    .B_N(_2091_),
    .Y(_2092_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5156_ (.Y(_2093_),
    .B(_2092_),
    .A_N(\falu_i.falutop.data_in[13] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5157_ (.A(\falu_i.falutop.data_in[14] ),
    .B(_1078_),
    .C(_2093_),
    .Y(_2094_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5158_ (.Y(_2095_),
    .B1(_2094_),
    .B2(net774),
    .A2(_1078_),
    .A1(net952),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5159_ (.VDD(VPWR),
    .Y(_0311_),
    .A(net953),
    .VSS(VGND));
 sg13g2_nor3_1 _5160_ (.A(\falu_i.falutop.data_in[0] ),
    .B(\falu_i.falutop.data_in[1] ),
    .C(\falu_i.falutop.data_in[2] ),
    .Y(_2096_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5161_ (.A(\falu_i.falutop.data_in[3] ),
    .B_N(_2096_),
    .Y(_2097_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5162_ (.A(\falu_i.falutop.data_in[4] ),
    .B_N(_2097_),
    .Y(_2098_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2b_1 _5163_ (.Y(_2099_),
    .B(_2098_),
    .A_N(\falu_i.falutop.data_in[5] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor3_1 _5164_ (.A(net1073),
    .B(net622),
    .C(_2099_),
    .Y(_2100_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a22oi_1 _5165_ (.Y(_2101_),
    .B1(net1074),
    .B2(net777),
    .A2(net622),
    .A1(net1054),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 _5166_ (.VDD(VPWR),
    .Y(_0312_),
    .A(net1075),
    .VSS(VGND));
 sg13g2_nor2_1 _5167_ (.A(net1148),
    .B(net620),
    .Y(_2102_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5168_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2301_),
    .A2(net620),
    .Y(_0313_),
    .B1(_2102_));
 sg13g2_nor2_1 _5169_ (.A(net1141),
    .B(net620),
    .Y(_2103_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5170_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2304_),
    .A2(net620),
    .Y(_0314_),
    .B1(_2103_));
 sg13g2_mux2_1 _5171_ (.A0(net1127),
    .A1(net765),
    .S(net618),
    .X(_0315_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5172_ (.A0(net1135),
    .A1(net760),
    .S(net618),
    .X(_0316_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5173_ (.A(net1114),
    .B(net617),
    .Y(_2104_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5174_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2303_),
    .A2(net617),
    .Y(_0317_),
    .B1(_2104_));
 sg13g2_nor2_1 _5175_ (.A(net1153),
    .B(net619),
    .Y(_2105_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5176_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2305_),
    .A2(net619),
    .Y(_0318_),
    .B1(_2105_));
 sg13g2_mux2_1 _5177_ (.A0(net1073),
    .A1(net749),
    .S(net618),
    .X(_0319_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5178_ (.A(net1137),
    .B(net619),
    .Y(_2106_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5179_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net705),
    .A2(net619),
    .Y(_0320_),
    .B1(_2106_));
 sg13g2_mux2_1 _5180_ (.A0(net1158),
    .A1(net743),
    .S(net618),
    .X(_0321_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5181_ (.A(net1123),
    .B(net618),
    .Y(_2107_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5182_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net707),
    .A2(net618),
    .Y(_0322_),
    .B1(_2107_));
 sg13g2_mux2_1 _5183_ (.A0(net1122),
    .A1(net735),
    .S(net618),
    .X(_0323_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5184_ (.A0(net1101),
    .A1(net730),
    .S(net618),
    .X(_0324_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5185_ (.A0(net1103),
    .A1(net725),
    .S(net617),
    .X(_0325_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5186_ (.A(net1086),
    .B(net617),
    .Y(_2108_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5187_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2296_),
    .A2(net617),
    .Y(_0326_),
    .B1(_2108_));
 sg13g2_nor2_1 _5188_ (.A(net1105),
    .B(net617),
    .Y(_2109_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5189_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(_2297_),
    .A2(net617),
    .Y(_0327_),
    .B1(_2109_));
 sg13g2_mux2_1 _5190_ (.A0(net776),
    .A1(net710),
    .S(net617),
    .X(_0328_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_mux2_1 _5191_ (.A0(net1081),
    .A1(\falu_i.falutop.data_in[0] ),
    .S(net624),
    .X(_0329_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5192_ (.Y(_2110_),
    .A(net413),
    .B(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5193_ (.Y(_2111_),
    .A(net777),
    .B(\falu_i.falutop.data_in[0] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5194_ (.B(_2111_),
    .A(\falu_i.falutop.data_in[1] ),
    .X(_2112_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5195_ (.B1(_2110_),
    .VDD(VPWR),
    .Y(_0330_),
    .VSS(VGND),
    .A1(net622),
    .A2(_2112_));
 sg13g2_nor2_1 _5196_ (.A(net891),
    .B(net624),
    .Y(_2113_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5197_ (.B1(net777),
    .VDD(VPWR),
    .Y(_2114_),
    .VSS(VGND),
    .A1(\falu_i.falutop.data_in[0] ),
    .A2(\falu_i.falutop.data_in[1] ));
 sg13g2_xor2_1 _5198_ (.B(_2114_),
    .A(\falu_i.falutop.data_in[2] ),
    .X(_2115_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5199_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net624),
    .A2(_2115_),
    .Y(_0331_),
    .B1(_2113_));
 sg13g2_nor2_1 _5200_ (.A(net967),
    .B(net623),
    .Y(_2116_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5201_ (.A(_2096_),
    .B_N(net777),
    .Y(_2117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5202_ (.Y(_2118_),
    .A(\falu_i.falutop.data_in[3] ),
    .B(_2117_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5203_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net623),
    .A2(_2118_),
    .Y(_0332_),
    .B1(_2116_));
 sg13g2_nor2_1 _5204_ (.A(net999),
    .B(net623),
    .Y(_2119_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5205_ (.A(_2097_),
    .B_N(net777),
    .Y(_2120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5206_ (.Y(_2121_),
    .A(\falu_i.falutop.data_in[4] ),
    .B(_2120_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5207_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net623),
    .A2(_2121_),
    .Y(_0333_),
    .B1(_2119_));
 sg13g2_nor2b_1 _5208_ (.A(_2098_),
    .B_N(net777),
    .Y(_2122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5209_ (.A(net983),
    .B(net623),
    .Y(_2123_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5210_ (.Y(_2124_),
    .A(\falu_i.falutop.data_in[5] ),
    .B(_2122_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5211_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net623),
    .A2(_2124_),
    .Y(_0334_),
    .B1(_2123_));
 sg13g2_nand2_1 _5212_ (.Y(_2125_),
    .A(net777),
    .B(_2099_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5213_ (.A(net920),
    .B(net623),
    .Y(_2126_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5214_ (.B(_2125_),
    .A(\falu_i.falutop.data_in[6] ),
    .X(_2127_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5215_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net623),
    .A2(_2127_),
    .Y(_0335_),
    .B1(_2126_));
 sg13g2_mux2_1 _5216_ (.A0(\falu_i.falutop.data_in[8] ),
    .A1(net906),
    .S(net622),
    .X(_0336_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5217_ (.Y(_2128_),
    .A(net388),
    .B(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5218_ (.Y(_2129_),
    .A(net775),
    .B(\falu_i.falutop.data_in[8] ),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5219_ (.B(_2129_),
    .A(\falu_i.falutop.data_in[9] ),
    .X(_2130_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5220_ (.B1(_2128_),
    .VDD(VPWR),
    .Y(_0337_),
    .VSS(VGND),
    .A1(net622),
    .A2(_2130_));
 sg13g2_nor2_1 _5221_ (.A(net475),
    .B(net625),
    .Y(_2131_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_o21ai_1 _5222_ (.B1(net776),
    .VDD(VPWR),
    .Y(_2132_),
    .VSS(VGND),
    .A1(\falu_i.falutop.data_in[8] ),
    .A2(\falu_i.falutop.data_in[9] ));
 sg13g2_xor2_1 _5223_ (.B(_2132_),
    .A(\falu_i.falutop.data_in[10] ),
    .X(_2133_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5224_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net625),
    .A2(_2133_),
    .Y(_0338_),
    .B1(_2131_));
 sg13g2_nor2b_1 _5225_ (.A(_2090_),
    .B_N(net776),
    .Y(_2134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5226_ (.A(net487),
    .B(net625),
    .Y(_2135_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5227_ (.Y(_2136_),
    .A(\falu_i.falutop.data_in[11] ),
    .B(_2134_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5228_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net625),
    .A2(_2136_),
    .Y(_0339_),
    .B1(_2135_));
 sg13g2_nor2_1 _5229_ (.A(net452),
    .B(net625),
    .Y(_2137_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2b_1 _5230_ (.A(_2091_),
    .B_N(net776),
    .Y(_2138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5231_ (.Y(_2139_),
    .A(\falu_i.falutop.data_in[12] ),
    .B(_2138_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5232_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net625),
    .A2(_2139_),
    .Y(_0340_),
    .B1(_2137_));
 sg13g2_nor2b_1 _5233_ (.A(_2092_),
    .B_N(net775),
    .Y(_2140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nor2_1 _5234_ (.A(net465),
    .B(net626),
    .Y(_2141_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xnor2_1 _5235_ (.Y(_2142_),
    .A(\falu_i.falutop.data_in[13] ),
    .B(_2140_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5236_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net626),
    .A2(_2142_),
    .Y(_0341_),
    .B1(_2141_));
 sg13g2_nor2_1 _5237_ (.A(net439),
    .B(net625),
    .Y(_2143_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_nand2_1 _5238_ (.Y(_2144_),
    .A(net773),
    .B(_2093_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_xor2_1 _5239_ (.B(_2144_),
    .A(\falu_i.falutop.data_in[14] ),
    .X(_2145_),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_a21oi_1 _5240_ (.VSS(VGND),
    .VDD(VPWR),
    .A1(net625),
    .A2(_2145_),
    .Y(_0342_),
    .B1(_2143_));
 sg13g2_dfrbpq_1 _5241_ (.RESET_B(net93),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0003_),
    .Q(\falu_i.falutop.i2c_inst.data_in[19] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5242_ (.RESET_B(net211),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0004_),
    .Q(\falu_i.falutop.i2c_inst.data_in[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5243_ (.RESET_B(net209),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0005_),
    .Q(\falu_i.falutop.i2c_inst.data_in[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5244_ (.RESET_B(net207),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0006_),
    .Q(\falu_i.falutop.i2c_inst.data_in[2] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5245_ (.RESET_B(net205),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0007_),
    .Q(\falu_i.falutop.i2c_inst.data_in[3] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_1 _5246_ (.RESET_B(net203),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0008_),
    .Q(\falu_i.falutop.i2c_inst.data_in[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5247_ (.RESET_B(net201),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0009_),
    .Q(\falu_i.falutop.i2c_inst.data_in[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5248_ (.RESET_B(net199),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0010_),
    .Q(\falu_i.falutop.i2c_inst.data_in[6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5249_ (.RESET_B(net197),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0011_),
    .Q(\falu_i.falutop.i2c_inst.data_in[7] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5250_ (.RESET_B(net195),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0012_),
    .Q(\falu_i.falutop.i2c_inst.data_in[8] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_1 _5251_ (.RESET_B(net193),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0013_),
    .Q(\falu_i.falutop.i2c_inst.data_in[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5252_ (.RESET_B(net191),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0014_),
    .Q(\falu_i.falutop.i2c_inst.data_in[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5253_ (.RESET_B(net189),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0015_),
    .Q(\falu_i.falutop.i2c_inst.data_in[11] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5254_ (.RESET_B(net187),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0016_),
    .Q(\falu_i.falutop.i2c_inst.data_in[12] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5255_ (.RESET_B(net185),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0017_),
    .Q(\falu_i.falutop.i2c_inst.data_in[13] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5256_ (.RESET_B(net183),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0018_),
    .Q(\falu_i.falutop.i2c_inst.data_in[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5257_ (.RESET_B(net181),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0019_),
    .Q(\falu_i.falutop.i2c_inst.data_in[15] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5258_ (.RESET_B(net179),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0020_),
    .Q(\falu_i.falutop.i2c_inst.data_in[16] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_1 _5259_ (.RESET_B(net177),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0021_),
    .Q(\falu_i.falutop.i2c_inst.data_in[17] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5260_ (.RESET_B(net175),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0022_),
    .Q(\falu_i.falutop.i2c_inst.data_in[18] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5261_ (.RESET_B(net173),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0023_),
    .Q(\ppwm_i.u_ppwm.u_mem.data_sync2 ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5262_ (.RESET_B(net172),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net382),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5263_ (.RESET_B(net170),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net507),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5264_ (.RESET_B(net168),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net521),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_1 _5265_ (.RESET_B(net166),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net458),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5266_ (.RESET_B(net164),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net471),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5267_ (.RESET_B(net162),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net427),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5268_ (.RESET_B(net160),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net493),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5269_ (.RESET_B(net158),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net431),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5270_ (.RESET_B(net156),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net925),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5271_ (.RESET_B(net154),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net536),
    .Q(\ppwm_i.u_ppwm.u_pwm.cmp_value[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _5272_ (.RESET_B(net152),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1113),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5273_ (.RESET_B(net150),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0035_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5274_ (.RESET_B(net148),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0036_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5275_ (.RESET_B(net146),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0037_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _5276_ (.RESET_B(net144),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1091),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _5277_ (.RESET_B(net142),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1061),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[5] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_1 _5278_ (.RESET_B(net140),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1068),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _5279_ (.RESET_B(net138),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0041_),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .CLK(clknet_leaf_14_clk));
 sg13g2_dfrbpq_2 _5280_ (.RESET_B(net136),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1095),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5281_ (.RESET_B(net134),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1025),
    .Q(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _5282_ (.RESET_B(net132),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net865),
    .Q(\ppwm_i.u_ppwm.period_start ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5283_ (.RESET_B(net131),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0045_),
    .Q(\ppwm_i.u_ppwm.global_counter[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5284_ (.RESET_B(net129),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net944),
    .Q(\ppwm_i.u_ppwm.global_counter[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5285_ (.RESET_B(net127),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1004),
    .Q(\ppwm_i.u_ppwm.global_counter[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_1 _5286_ (.RESET_B(net125),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0048_),
    .Q(\ppwm_i.u_ppwm.global_counter[3] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5287_ (.RESET_B(net123),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1109),
    .Q(\ppwm_i.u_ppwm.global_counter[4] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5288_ (.RESET_B(net121),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1147),
    .Q(\ppwm_i.u_ppwm.global_counter[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_1 _5289_ (.RESET_B(net119),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0051_),
    .Q(\ppwm_i.u_ppwm.global_counter[6] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5290_ (.RESET_B(net117),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0052_),
    .Q(\ppwm_i.u_ppwm.global_counter[7] ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _5291_ (.RESET_B(net115),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net555),
    .Q(\ppwm_i.u_ppwm.global_counter[8] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5292_ (.RESET_B(net113),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0054_),
    .Q(\ppwm_i.u_ppwm.global_counter[9] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5293_ (.RESET_B(net111),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0055_),
    .Q(\ppwm_i.u_ppwm.global_counter[10] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5294_ (.RESET_B(net109),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net956),
    .Q(\ppwm_i.u_ppwm.global_counter[11] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5295_ (.RESET_B(net107),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0057_),
    .Q(\ppwm_i.u_ppwm.global_counter[12] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5296_ (.RESET_B(net105),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0058_),
    .Q(\ppwm_i.u_ppwm.global_counter[13] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5297_ (.RESET_B(net103),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net976),
    .Q(\ppwm_i.u_ppwm.global_counter[14] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5298_ (.RESET_B(net101),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0060_),
    .Q(\ppwm_i.u_ppwm.global_counter[15] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5299_ (.RESET_B(net99),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0061_),
    .Q(\ppwm_i.u_ppwm.global_counter[16] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5300_ (.RESET_B(net97),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net991),
    .Q(\ppwm_i.u_ppwm.global_counter[17] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5301_ (.RESET_B(net92),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1077),
    .Q(\ppwm_i.u_ppwm.global_counter[18] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5302_ (.RESET_B(net90),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1032),
    .Q(\ppwm_i.u_ppwm.global_counter[19] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_1 _5303_ (.RESET_B(net94),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net377),
    .Q(\ppwm_i.u_ppwm.data_o ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_1 _5304_ (.RESET_B(net95),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net982),
    .Q(\ppwm_i.u_ppwm.u_ex.state_q[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5305_ (.RESET_B(net223),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net387),
    .Q(\ppwm_i.u_ppwm.u_ex.state_q[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5306_ (.RESET_B(net88),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1040),
    .Q(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _5307_ (.RESET_B(net87),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1164),
    .Q(\ppwm_i.u_ppwm.pc[0] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5308_ (.RESET_B(net85),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0067_),
    .Q(\ppwm_i.u_ppwm.pc[1] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5309_ (.RESET_B(net83),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0068_),
    .Q(\ppwm_i.u_ppwm.pc[2] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5310_ (.RESET_B(net81),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0069_),
    .Q(\ppwm_i.u_ppwm.pc[3] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_2 _5311_ (.RESET_B(net79),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0070_),
    .Q(\ppwm_i.u_ppwm.u_ex.cmp_flag_q ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _5312_ (.RESET_B(net77),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0071_),
    .Q(\ppwm_i.u_ppwm.polarity ),
    .CLK(clknet_leaf_15_clk));
 sg13g2_dfrbpq_2 _5313_ (.RESET_B(net75),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0072_),
    .Q(\ppwm_i.u_ppwm.pwm_value[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5314_ (.RESET_B(net73),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1197),
    .Q(\ppwm_i.u_ppwm.pwm_value[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5315_ (.RESET_B(net71),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0074_),
    .Q(\ppwm_i.u_ppwm.pwm_value[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5316_ (.RESET_B(net69),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0075_),
    .Q(\ppwm_i.u_ppwm.pwm_value[3] ),
    .CLK(clknet_leaf_12_clk));
 sg13g2_dfrbpq_2 _5317_ (.RESET_B(net67),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1182),
    .Q(\ppwm_i.u_ppwm.pwm_value[4] ),
    .CLK(clknet_leaf_18_clk));
 sg13g2_dfrbpq_2 _5318_ (.RESET_B(net65),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0077_),
    .Q(\ppwm_i.u_ppwm.pwm_value[5] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5319_ (.RESET_B(net63),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0078_),
    .Q(\ppwm_i.u_ppwm.pwm_value[6] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5320_ (.RESET_B(net61),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1191),
    .Q(\ppwm_i.u_ppwm.pwm_value[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5321_ (.RESET_B(net59),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0080_),
    .Q(\ppwm_i.u_ppwm.pwm_value[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5322_ (.RESET_B(net57),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0081_),
    .Q(\ppwm_i.u_ppwm.pwm_value[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5323_ (.RESET_B(net55),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0082_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_2 _5324_ (.RESET_B(net53),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0083_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5325_ (.RESET_B(net51),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0084_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5326_ (.RESET_B(net49),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0085_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5327_ (.RESET_B(net47),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0086_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .CLK(clknet_leaf_13_clk));
 sg13g2_dfrbpq_2 _5328_ (.RESET_B(net45),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1175),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .CLK(clknet_leaf_16_clk));
 sg13g2_dfrbpq_2 _5329_ (.RESET_B(net43),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0088_),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5330_ (.RESET_B(net41),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1170),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _5331_ (.RESET_B(net39),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1195),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_2 _5332_ (.RESET_B(net37),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1161),
    .Q(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .CLK(clknet_leaf_17_clk));
 sg13g2_dfrbpq_1 _5333_ (.RESET_B(net35),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net421),
    .Q(\falu_i.falutop.i2c_inst.op[0] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5334_ (.RESET_B(net34),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net913),
    .Q(\falu_i.falutop.i2c_inst.op[1] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5335_ (.RESET_B(net33),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net468),
    .Q(\falu_i.falutop.i2c_inst.op[2] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5336_ (.RESET_B(net32),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net429),
    .Q(\falu_i.falutop.i2c_inst.op[3] ),
    .CLK(clknet_leaf_19_clk));
 sg13g2_dfrbpq_1 _5337_ (.RESET_B(net31),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0096_),
    .Q(\ppwm_i.u_ppwm.u_mem.clk_prog_sync1 ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5338_ (.RESET_B(net30),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0097_),
    .Q(\ppwm_i.u_ppwm.u_mem.clk_prog_sync2 ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5339_ (.RESET_B(net372),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0098_),
    .Q(\ppwm_i.u_ppwm.u_mem.clk_prog_sync3 ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5340_ (.RESET_B(net371),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0099_),
    .Q(\ppwm_i.u_ppwm.u_mem.data_sync1 ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_1 _5341_ (.RESET_B(net370),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0100_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[0] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5342_ (.RESET_B(net368),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net524),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[1] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5343_ (.RESET_B(net366),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net853),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[2] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5344_ (.RESET_B(net364),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net561),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[3] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5345_ (.RESET_B(net362),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0104_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[4] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5346_ (.RESET_B(net360),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net484),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5347_ (.RESET_B(net358),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0106_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[6] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5348_ (.RESET_B(net356),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0107_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[7] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5349_ (.RESET_B(net354),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net442),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[8] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5350_ (.RESET_B(net352),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net505),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[9] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5351_ (.RESET_B(net350),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0110_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[10] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5352_ (.RESET_B(net348),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0111_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[11] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5353_ (.RESET_B(net346),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0112_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[12] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5354_ (.RESET_B(net344),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net929),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5355_ (.RESET_B(net342),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net497),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[14] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5356_ (.RESET_B(net340),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0115_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[15] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5357_ (.RESET_B(net338),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net448),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5358_ (.RESET_B(net336),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0117_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[17] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5359_ (.RESET_B(net334),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0118_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[18] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5360_ (.RESET_B(net332),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net876),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[19] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_2 _5361_ (.RESET_B(net330),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net966),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[20] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5362_ (.RESET_B(net328),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net478),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[21] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5363_ (.RESET_B(net326),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0122_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[22] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5364_ (.RESET_B(net324),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net403),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .CLK(clknet_leaf_33_clk));
 sg13g2_dfrbpq_1 _5365_ (.RESET_B(net322),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0124_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[24] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5366_ (.RESET_B(net320),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net509),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[25] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5367_ (.RESET_B(net318),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0126_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[26] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_1 _5368_ (.RESET_B(net316),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net960),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5369_ (.RESET_B(net314),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0128_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[28] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5370_ (.RESET_B(net312),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net846),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[29] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5371_ (.RESET_B(net310),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net517),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[30] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5372_ (.RESET_B(net308),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0131_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[31] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5373_ (.RESET_B(net306),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0132_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[32] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5374_ (.RESET_B(net304),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net548),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[33] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5375_ (.RESET_B(net302),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0134_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5376_ (.RESET_B(net300),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net473),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[35] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5377_ (.RESET_B(net298),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0136_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[36] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5378_ (.RESET_B(net296),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net425),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[37] ),
    .CLK(clknet_leaf_21_clk));
 sg13g2_dfrbpq_1 _5379_ (.RESET_B(net294),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net423),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[38] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5380_ (.RESET_B(net292),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0139_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[39] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5381_ (.RESET_B(net290),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net456),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[40] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5382_ (.RESET_B(net288),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net970),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[41] ),
    .CLK(clknet_leaf_22_clk));
 sg13g2_dfrbpq_1 _5383_ (.RESET_B(net286),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net855),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[42] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5384_ (.RESET_B(net284),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0143_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[43] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5385_ (.RESET_B(net282),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0144_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[44] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5386_ (.RESET_B(net280),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net531),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[45] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5387_ (.RESET_B(net278),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0146_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[46] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5388_ (.RESET_B(net276),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0147_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[47] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_2 _5389_ (.RESET_B(net274),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0148_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[48] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5390_ (.RESET_B(net272),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0149_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[49] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5391_ (.RESET_B(net270),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net408),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[50] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5392_ (.RESET_B(net268),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net916),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[51] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5393_ (.RESET_B(net266),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net444),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[52] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_1 _5394_ (.RESET_B(net264),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0153_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[53] ),
    .CLK(clknet_leaf_23_clk));
 sg13g2_dfrbpq_1 _5395_ (.RESET_B(net262),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0154_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[54] ),
    .CLK(clknet_leaf_24_clk));
 sg13g2_dfrbpq_2 _5396_ (.RESET_B(net260),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0155_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[55] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5397_ (.RESET_B(net258),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net395),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[56] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5398_ (.RESET_B(net256),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net558),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[57] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5399_ (.RESET_B(net254),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0158_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[58] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5400_ (.RESET_B(net252),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0159_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[59] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5401_ (.RESET_B(net250),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net438),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[60] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5402_ (.RESET_B(net248),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0161_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[61] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _5403_ (.RESET_B(net246),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0162_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[62] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5404_ (.RESET_B(net244),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net450),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[63] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5405_ (.RESET_B(net242),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0164_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[64] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5406_ (.RESET_B(net240),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0165_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[65] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5407_ (.RESET_B(net238),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net890),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[66] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5408_ (.RESET_B(net236),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0167_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[67] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5409_ (.RESET_B(net234),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0168_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[68] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5410_ (.RESET_B(net232),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net464),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5411_ (.RESET_B(net230),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net416),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[70] ),
    .CLK(clknet_leaf_25_clk));
 sg13g2_dfrbpq_1 _5412_ (.RESET_B(net228),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0171_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[71] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5413_ (.RESET_B(net226),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0172_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[72] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5414_ (.RESET_B(net224),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net923),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[73] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5415_ (.RESET_B(net222),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net384),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[74] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5416_ (.RESET_B(net220),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0175_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[75] ),
    .CLK(clknet_leaf_27_clk));
 sg13g2_dfrbpq_1 _5417_ (.RESET_B(net218),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0176_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[76] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5418_ (.RESET_B(net216),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net552),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[77] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5419_ (.RESET_B(net214),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net546),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[78] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_1 _5420_ (.RESET_B(net212),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0179_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[79] ),
    .CLK(clknet_leaf_26_clk));
 sg13g2_dfrbpq_2 _5421_ (.RESET_B(net208),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0180_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[80] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _5422_ (.RESET_B(net204),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net418),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[81] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _5423_ (.RESET_B(net200),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0182_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[82] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5424_ (.RESET_B(net196),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0183_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[83] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _5425_ (.RESET_B(net192),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0184_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[84] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5426_ (.RESET_B(net188),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net511),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[85] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5427_ (.RESET_B(net184),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0186_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5428_ (.RESET_B(net180),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net519),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[87] ),
    .CLK(clknet_leaf_29_clk));
 sg13g2_dfrbpq_1 _5429_ (.RESET_B(net176),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0188_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5430_ (.RESET_B(net171),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net503),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[89] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5431_ (.RESET_B(net167),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net958),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[90] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5432_ (.RESET_B(net163),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net391),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[91] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5433_ (.RESET_B(net159),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0192_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[92] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5434_ (.RESET_B(net155),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0193_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[93] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5435_ (.RESET_B(net151),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0194_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[94] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _5436_ (.RESET_B(net147),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0195_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[95] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_1 _5437_ (.RESET_B(net143),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net533),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[96] ),
    .CLK(clknet_leaf_28_clk));
 sg13g2_dfrbpq_2 _5438_ (.RESET_B(net139),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0197_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5439_ (.RESET_B(net135),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0198_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[98] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5440_ (.RESET_B(net130),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net538),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[99] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_2 _5441_ (.RESET_B(net126),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net501),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[100] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5442_ (.RESET_B(net122),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0201_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[101] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5443_ (.RESET_B(net118),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net393),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[102] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5444_ (.RESET_B(net114),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0203_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[103] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_2 _5445_ (.RESET_B(net110),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0204_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[104] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5446_ (.RESET_B(net106),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net529),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[105] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5447_ (.RESET_B(net102),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net446),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[106] ),
    .CLK(clknet_leaf_30_clk));
 sg13g2_dfrbpq_1 _5448_ (.RESET_B(net98),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0207_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[107] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5449_ (.RESET_B(net91),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net462),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[108] ),
    .CLK(clknet_leaf_31_clk));
 sg13g2_dfrbpq_1 _5450_ (.RESET_B(net86),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0209_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[109] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5451_ (.RESET_B(net82),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0210_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[110] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_1 _5452_ (.RESET_B(net78),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0211_),
    .Q(\ppwm_i.u_ppwm.u_mem.memory[111] ),
    .CLK(clknet_leaf_32_clk));
 sg13g2_dfrbpq_2 _5453_ (.RESET_B(net74),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net379),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[0] ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5454_ (.RESET_B(net70),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0213_),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[1] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5455_ (.RESET_B(net66),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1053),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[2] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5456_ (.RESET_B(net62),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0215_),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _5457_ (.RESET_B(net58),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1012),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _5458_ (.RESET_B(net54),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1157),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_1 _5459_ (.RESET_B(net50),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net514),
    .Q(\ppwm_i.u_ppwm.u_mem.bit_count[6] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_2 _5460_ (.RESET_B(net46),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net936),
    .Q(\ppwm_i.u_ppwm.u_mem.programming ),
    .CLK(clknet_leaf_11_clk));
 sg13g2_dfrbpq_2 _5461_ (.RESET_B(net42),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net460),
    .Q(\falu_i.falutop.i2c_inst.state[0] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5462_ (.RESET_B(net38),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0221_),
    .Q(\falu_i.falutop.i2c_inst.state[1] ),
    .CLK(clknet_leaf_9_clk));
 sg13g2_dfrbpq_2 _5463_ (.RESET_B(net369),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0222_),
    .Q(\falu_i.falutop.i2c_inst.counter[0] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _5464_ (.RESET_B(net365),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0223_),
    .Q(\falu_i.falutop.i2c_inst.counter[1] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _5465_ (.RESET_B(net361),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0224_),
    .Q(\falu_i.falutop.i2c_inst.counter[2] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _5466_ (.RESET_B(net357),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0225_),
    .Q(\falu_i.falutop.i2c_inst.counter[3] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _5467_ (.RESET_B(net353),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0226_),
    .Q(\falu_i.falutop.i2c_inst.counter[4] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5468_ (.RESET_B(net349),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0227_),
    .Q(\falu_i.falutop.div_inst.start ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _5469_ (.RESET_B(net347),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net849),
    .Q(\falu_i.falutop.data_in[0] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5470_ (.RESET_B(net345),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net902),
    .Q(\falu_i.falutop.data_in[1] ),
    .CLK(clknet_leaf_8_clk));
 sg13g2_dfrbpq_2 _5471_ (.RESET_B(net343),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net973),
    .Q(\falu_i.falutop.data_in[2] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5472_ (.RESET_B(net341),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net993),
    .Q(\falu_i.falutop.data_in[3] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5473_ (.RESET_B(net339),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net882),
    .Q(\falu_i.falutop.data_in[4] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5474_ (.RESET_B(net337),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net870),
    .Q(\falu_i.falutop.data_in[5] ),
    .CLK(clknet_leaf_10_clk));
 sg13g2_dfrbpq_2 _5475_ (.RESET_B(net335),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net851),
    .Q(\falu_i.falutop.data_in[6] ),
    .CLK(clknet_leaf_5_clk));
 sg13g2_dfrbpq_2 _5476_ (.RESET_B(net333),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net872),
    .Q(\falu_i.falutop.data_in[7] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5477_ (.RESET_B(net331),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net874),
    .Q(\falu_i.falutop.data_in[8] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5478_ (.RESET_B(net329),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net900),
    .Q(\falu_i.falutop.data_in[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5479_ (.RESET_B(net327),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net946),
    .Q(\falu_i.falutop.data_in[10] ),
    .CLK(clknet_leaf_7_clk));
 sg13g2_dfrbpq_2 _5480_ (.RESET_B(net325),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net859),
    .Q(\falu_i.falutop.data_in[11] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5481_ (.RESET_B(net323),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net927),
    .Q(\falu_i.falutop.data_in[12] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5482_ (.RESET_B(net321),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net895),
    .Q(\falu_i.falutop.data_in[13] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5483_ (.RESET_B(net319),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net862),
    .Q(\falu_i.falutop.data_in[14] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5484_ (.RESET_B(net317),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net909),
    .Q(\falu_i.falutop.data_in[15] ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_1 _5485_ (.RESET_B(net315),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net998),
    .Q(\falu_i.falutop.i2c_inst.sda_o ),
    .CLK(clknet_leaf_6_clk));
 sg13g2_dfrbpq_2 _5486_ (.RESET_B(net311),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0245_),
    .Q(\falu_i.falutop.div_inst.acc[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _5487_ (.RESET_B(net309),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0246_),
    .Q(\falu_i.falutop.div_inst.quo[0] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5488_ (.RESET_B(net305),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0247_),
    .Q(\falu_i.falutop.div_inst.done ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5489_ (.RESET_B(net303),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0248_),
    .Q(\falu_i.falutop.alu_inst.op[0] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _5490_ (.RESET_B(net301),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0249_),
    .Q(\falu_i.falutop.alu_inst.op[1] ),
    .CLK(clknet_leaf_20_clk));
 sg13g2_dfrbpq_2 _5491_ (.RESET_B(net299),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0250_),
    .Q(\falu_i.falutop.alu_inst.op[2] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_2 _5492_ (.RESET_B(net297),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0251_),
    .Q(\falu_i.falutop.alu_inst.op[3] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _5493_ (.RESET_B(net295),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net527),
    .Q(\falu_i.falutop.div_inst.i[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _5494_ (.RESET_B(net291),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net919),
    .Q(\falu_i.falutop.div_inst.i[1] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _5495_ (.RESET_B(net287),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net410),
    .Q(\falu_i.falutop.div_inst.i[2] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _5496_ (.RESET_B(net283),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0255_),
    .Q(\falu_i.falutop.div_inst.b1[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5497_ (.RESET_B(net281),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0256_),
    .Q(\falu_i.falutop.div_inst.b1[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5498_ (.RESET_B(net279),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0257_),
    .Q(\falu_i.falutop.div_inst.b1[2] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5499_ (.RESET_B(net277),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0258_),
    .Q(\falu_i.falutop.div_inst.b1[3] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5500_ (.RESET_B(net275),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0259_),
    .Q(\falu_i.falutop.div_inst.b1[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5501_ (.RESET_B(net273),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0260_),
    .Q(\falu_i.falutop.div_inst.b1[5] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5502_ (.RESET_B(net271),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0261_),
    .Q(\falu_i.falutop.div_inst.b1[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_2 _5503_ (.RESET_B(net269),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1055),
    .Q(\falu_i.falutop.div_inst.b1[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5504_ (.RESET_B(net267),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0263_),
    .Q(\falu_i.falutop.div_inst.busy ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_2 _5505_ (.RESET_B(net265),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0264_),
    .Q(\falu_i.falutop.div_inst.val[0] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_2 _5506_ (.RESET_B(net261),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net941),
    .Q(\falu_i.falutop.div_inst.val[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _5507_ (.RESET_B(net257),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net979),
    .Q(\falu_i.falutop.div_inst.val[2] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5508_ (.RESET_B(net253),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0267_),
    .Q(\falu_i.falutop.div_inst.val[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5509_ (.RESET_B(net249),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0268_),
    .Q(\falu_i.falutop.div_inst.val[4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5510_ (.RESET_B(net245),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0269_),
    .Q(\falu_i.falutop.div_inst.val[5] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5511_ (.RESET_B(net241),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1038),
    .Q(\falu_i.falutop.div_inst.val[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _5512_ (.RESET_B(net237),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net543),
    .Q(\falu_i.falutop.div_inst.val[7] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_2 _5513_ (.RESET_B(net233),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0272_),
    .Q(\falu_i.falutop.div_inst.rem[0] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5514_ (.RESET_B(net229),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1099),
    .Q(\falu_i.falutop.div_inst.rem[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5515_ (.RESET_B(net225),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0274_),
    .Q(\falu_i.falutop.div_inst.rem[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5516_ (.RESET_B(net221),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0275_),
    .Q(\falu_i.falutop.div_inst.rem[3] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5517_ (.RESET_B(net217),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0276_),
    .Q(\falu_i.falutop.div_inst.rem[4] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_1 _5518_ (.RESET_B(net213),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0277_),
    .Q(\falu_i.falutop.div_inst.rem[5] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5519_ (.RESET_B(net206),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0278_),
    .Q(\falu_i.falutop.div_inst.rem[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5520_ (.RESET_B(net198),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0279_),
    .Q(\falu_i.falutop.div_inst.rem[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _5521_ (.RESET_B(net190),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net400),
    .Q(\falu_i.falutop.div_inst.quo[1] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _5522_ (.RESET_B(net186),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net412),
    .Q(\falu_i.falutop.div_inst.quo[2] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5523_ (.RESET_B(net182),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net436),
    .Q(\falu_i.falutop.div_inst.quo[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5524_ (.RESET_B(net178),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net406),
    .Q(\falu_i.falutop.div_inst.quo[4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5525_ (.RESET_B(net174),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net433),
    .Q(\falu_i.falutop.div_inst.quo[5] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5526_ (.RESET_B(net169),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0285_),
    .Q(\falu_i.falutop.div_inst.quo[6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _5527_ (.RESET_B(net165),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net397),
    .Q(\falu_i.falutop.div_inst.acc_next[0] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_2 _5528_ (.RESET_B(net161),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net499),
    .Q(\falu_i.falutop.div_inst.acc[1] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5529_ (.RESET_B(net153),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net490),
    .Q(\falu_i.falutop.div_inst.acc[2] ),
    .CLK(clknet_leaf_1_clk));
 sg13g2_dfrbpq_2 _5530_ (.RESET_B(net145),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net495),
    .Q(\falu_i.falutop.div_inst.acc[3] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5531_ (.RESET_B(net137),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net857),
    .Q(\falu_i.falutop.div_inst.acc[4] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5532_ (.RESET_B(net128),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net550),
    .Q(\falu_i.falutop.div_inst.acc[5] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_2 _5533_ (.RESET_B(net120),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net932),
    .Q(\falu_i.falutop.div_inst.acc[6] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5534_ (.RESET_B(net112),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net486),
    .Q(\falu_i.falutop.div_inst.acc[7] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5535_ (.RESET_B(net104),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0294_),
    .Q(\falu_i.falutop.div_inst.acc[8] ),
    .CLK(clknet_leaf_0_clk));
 sg13g2_dfrbpq_1 _5536_ (.RESET_B(net96),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1023),
    .Q(\falu_i.falutop.i2c_inst.result[0] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _5537_ (.RESET_B(net84),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1058),
    .Q(\falu_i.falutop.i2c_inst.result[1] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5538_ (.RESET_B(net76),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1048),
    .Q(\falu_i.falutop.i2c_inst.result[2] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _5539_ (.RESET_B(net68),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0298_),
    .Q(\falu_i.falutop.i2c_inst.result[3] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_1 _5540_ (.RESET_B(net60),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0299_),
    .Q(\falu_i.falutop.i2c_inst.result[4] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5541_ (.RESET_B(net52),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0300_),
    .Q(\falu_i.falutop.i2c_inst.result[5] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _5542_ (.RESET_B(net44),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0301_),
    .Q(\falu_i.falutop.i2c_inst.result[6] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _5543_ (.RESET_B(net36),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1042),
    .Q(\falu_i.falutop.i2c_inst.result[7] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5544_ (.RESET_B(net363),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1034),
    .Q(\falu_i.falutop.i2c_inst.result[8] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5545_ (.RESET_B(net355),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1065),
    .Q(\falu_i.falutop.i2c_inst.result[9] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5546_ (.RESET_B(net313),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1063),
    .Q(\falu_i.falutop.i2c_inst.result[10] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5547_ (.RESET_B(net293),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1021),
    .Q(\falu_i.falutop.i2c_inst.result[11] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5548_ (.RESET_B(net285),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1019),
    .Q(\falu_i.falutop.i2c_inst.result[12] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5549_ (.RESET_B(net259),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1036),
    .Q(\falu_i.falutop.i2c_inst.result[13] ),
    .CLK(clknet_leaf_39_clk));
 sg13g2_dfrbpq_1 _5550_ (.RESET_B(net251),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1072),
    .Q(\falu_i.falutop.i2c_inst.result[14] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5551_ (.RESET_B(net243),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1030),
    .Q(\falu_i.falutop.i2c_inst.result[15] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5552_ (.RESET_B(net235),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0311_),
    .Q(\falu_i.falutop.div_inst.a[7] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_dfrbpq_1 _5553_ (.RESET_B(net227),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0312_),
    .Q(\falu_i.falutop.div_inst.b[7] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5554_ (.RESET_B(net219),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1149),
    .Q(\falu_i.falutop.alu_data_in[0] ),
    .CLK(clknet_leaf_34_clk));
 sg13g2_dfrbpq_1 _5555_ (.RESET_B(net215),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1142),
    .Q(\falu_i.falutop.alu_data_in[1] ),
    .CLK(clknet_leaf_35_clk));
 sg13g2_dfrbpq_1 _5556_ (.RESET_B(net210),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1128),
    .Q(\falu_i.falutop.alu_data_in[2] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5557_ (.RESET_B(net202),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1136),
    .Q(\falu_i.falutop.alu_data_in[3] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5558_ (.RESET_B(net194),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1115),
    .Q(\falu_i.falutop.alu_data_in[4] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5559_ (.RESET_B(net157),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1154),
    .Q(\falu_i.falutop.alu_data_in[5] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _5560_ (.RESET_B(net149),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0319_),
    .Q(\falu_i.falutop.alu_data_in[6] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5561_ (.RESET_B(net141),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1138),
    .Q(\falu_i.falutop.alu_data_in[7] ),
    .CLK(clknet_leaf_36_clk));
 sg13g2_dfrbpq_1 _5562_ (.RESET_B(net133),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1159),
    .Q(\falu_i.falutop.alu_data_in[8] ),
    .CLK(clknet_leaf_38_clk));
 sg13g2_dfrbpq_2 _5563_ (.RESET_B(net124),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0322_),
    .Q(\falu_i.falutop.alu_data_in[9] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_1 _5564_ (.RESET_B(net116),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0323_),
    .Q(\falu_i.falutop.alu_data_in[10] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5565_ (.RESET_B(net108),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1102),
    .Q(\falu_i.falutop.alu_data_in[11] ),
    .CLK(clknet_leaf_37_clk));
 sg13g2_dfrbpq_2 _5566_ (.RESET_B(net100),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1104),
    .Q(\falu_i.falutop.alu_data_in[12] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_2 _5567_ (.RESET_B(net89),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1087),
    .Q(\falu_i.falutop.alu_data_in[13] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _5568_ (.RESET_B(net80),
    .VSS(VGND),
    .VDD(VPWR),
    .D(_0327_),
    .Q(\falu_i.falutop.alu_data_in[14] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _5569_ (.RESET_B(net72),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1179),
    .Q(\falu_i.falutop.alu_data_in[15] ),
    .CLK(clknet_leaf_40_clk));
 sg13g2_dfrbpq_1 _5570_ (.RESET_B(net64),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1082),
    .Q(\falu_i.falutop.div_inst.b[0] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5571_ (.RESET_B(net56),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net414),
    .Q(\falu_i.falutop.div_inst.b[1] ),
    .CLK(clknet_leaf_2_clk));
 sg13g2_dfrbpq_1 _5572_ (.RESET_B(net48),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net892),
    .Q(\falu_i.falutop.div_inst.b[2] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5573_ (.RESET_B(net40),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net968),
    .Q(\falu_i.falutop.div_inst.b[3] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5574_ (.RESET_B(net367),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net1000),
    .Q(\falu_i.falutop.div_inst.b[4] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5575_ (.RESET_B(net359),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net984),
    .Q(\falu_i.falutop.div_inst.b[5] ),
    .CLK(clknet_leaf_4_clk));
 sg13g2_dfrbpq_1 _5576_ (.RESET_B(net351),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net921),
    .Q(\falu_i.falutop.div_inst.b[6] ),
    .CLK(clknet_leaf_3_clk));
 sg13g2_dfrbpq_1 _5577_ (.RESET_B(net307),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net907),
    .Q(\falu_i.falutop.div_inst.a[0] ),
    .CLK(clknet_leaf_44_clk));
 sg13g2_dfrbpq_1 _5578_ (.RESET_B(net289),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net389),
    .Q(\falu_i.falutop.div_inst.a[1] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5579_ (.RESET_B(net263),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net476),
    .Q(\falu_i.falutop.div_inst.a[2] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5580_ (.RESET_B(net255),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net488),
    .Q(\falu_i.falutop.div_inst.a[3] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5581_ (.RESET_B(net247),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net453),
    .Q(\falu_i.falutop.div_inst.a[4] ),
    .CLK(clknet_leaf_41_clk));
 sg13g2_dfrbpq_1 _5582_ (.RESET_B(net239),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net466),
    .Q(\falu_i.falutop.div_inst.a[5] ),
    .CLK(clknet_leaf_42_clk));
 sg13g2_dfrbpq_1 _5583_ (.RESET_B(net231),
    .VSS(VGND),
    .VDD(VPWR),
    .D(net440),
    .Q(\falu_i.falutop.div_inst.a[6] ),
    .CLK(clknet_leaf_43_clk));
 sg13g2_tiehi _5337__31 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net31));
 sg13g2_tiehi _5336__32 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net32));
 sg13g2_tiehi _5335__33 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net33));
 sg13g2_tiehi _5334__34 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net34));
 sg13g2_tiehi _5333__35 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net35));
 sg13g2_tiehi _5543__36 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net36));
 sg13g2_tiehi _5332__37 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net37));
 sg13g2_tiehi _5462__38 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net38));
 sg13g2_tiehi _5331__39 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net39));
 sg13g2_tiehi _5573__40 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net40));
 sg13g2_tiehi _5330__41 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net41));
 sg13g2_tiehi _5461__42 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net42));
 sg13g2_tiehi _5329__43 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net43));
 sg13g2_tiehi _5542__44 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net44));
 sg13g2_tiehi _5328__45 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net45));
 sg13g2_tiehi _5460__46 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net46));
 sg13g2_tiehi _5327__47 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net47));
 sg13g2_tiehi _5572__48 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net48));
 sg13g2_tiehi _5326__49 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net49));
 sg13g2_tiehi _5459__50 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net50));
 sg13g2_tiehi _5325__51 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net51));
 sg13g2_tiehi _5541__52 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net52));
 sg13g2_tiehi _5324__53 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net53));
 sg13g2_tiehi _5458__54 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net54));
 sg13g2_tiehi _5323__55 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net55));
 sg13g2_tiehi _5571__56 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net56));
 sg13g2_tiehi _5322__57 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net57));
 sg13g2_tiehi _5457__58 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net58));
 sg13g2_tiehi _5321__59 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net59));
 sg13g2_tiehi _5540__60 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net60));
 sg13g2_tiehi _5320__61 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net61));
 sg13g2_tiehi _5456__62 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net62));
 sg13g2_tiehi _5319__63 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net63));
 sg13g2_tiehi _5570__64 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net64));
 sg13g2_tiehi _5318__65 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net65));
 sg13g2_tiehi _5455__66 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net66));
 sg13g2_tiehi _5317__67 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net67));
 sg13g2_tiehi _5539__68 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net68));
 sg13g2_tiehi _5316__69 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net69));
 sg13g2_tiehi _5454__70 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net70));
 sg13g2_tiehi _5315__71 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net71));
 sg13g2_tiehi _5569__72 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net72));
 sg13g2_tiehi _5314__73 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net73));
 sg13g2_tiehi _5453__74 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net74));
 sg13g2_tiehi _5313__75 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net75));
 sg13g2_tiehi _5538__76 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net76));
 sg13g2_tiehi _5312__77 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net77));
 sg13g2_tiehi _5452__78 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net78));
 sg13g2_tiehi _5311__79 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net79));
 sg13g2_tiehi _5568__80 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net80));
 sg13g2_tiehi _5310__81 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net81));
 sg13g2_tiehi _5451__82 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net82));
 sg13g2_tiehi _5309__83 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net83));
 sg13g2_tiehi _5537__84 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net84));
 sg13g2_tiehi _5308__85 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net85));
 sg13g2_tiehi _5450__86 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net86));
 sg13g2_tiehi _5307__87 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net87));
 sg13g2_tiehi _5306__88 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net88));
 sg13g2_tiehi _5567__89 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net89));
 sg13g2_tiehi _5302__90 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net90));
 sg13g2_tiehi _5449__91 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net91));
 sg13g2_tiehi _5301__92 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net92));
 sg13g2_tiehi _5241__93 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net93));
 sg13g2_tiehi _5303__94 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net94));
 sg13g2_tiehi _5304__95 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net95));
 sg13g2_tiehi _5536__96 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net96));
 sg13g2_tiehi _5300__97 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net97));
 sg13g2_tiehi _5448__98 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net98));
 sg13g2_tiehi _5299__99 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net99));
 sg13g2_tiehi _5566__100 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net100));
 sg13g2_tiehi _5298__101 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net101));
 sg13g2_tiehi _5447__102 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net102));
 sg13g2_tiehi _5297__103 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net103));
 sg13g2_tiehi _5535__104 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net104));
 sg13g2_tiehi _5296__105 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net105));
 sg13g2_tiehi _5446__106 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net106));
 sg13g2_tiehi _5295__107 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net107));
 sg13g2_tiehi _5565__108 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net108));
 sg13g2_tiehi _5294__109 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net109));
 sg13g2_tiehi _5445__110 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net110));
 sg13g2_tiehi _5293__111 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net111));
 sg13g2_tiehi _5534__112 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net112));
 sg13g2_tiehi _5292__113 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net113));
 sg13g2_tiehi _5444__114 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net114));
 sg13g2_tiehi _5291__115 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net115));
 sg13g2_tiehi _5564__116 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net116));
 sg13g2_tiehi _5290__117 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net117));
 sg13g2_tiehi _5443__118 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net118));
 sg13g2_tiehi _5289__119 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net119));
 sg13g2_tiehi _5533__120 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net120));
 sg13g2_tiehi _5288__121 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net121));
 sg13g2_tiehi _5442__122 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net122));
 sg13g2_tiehi _5287__123 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net123));
 sg13g2_tiehi _5563__124 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net124));
 sg13g2_tiehi _5286__125 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net125));
 sg13g2_tiehi _5441__126 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net126));
 sg13g2_tiehi _5285__127 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net127));
 sg13g2_tiehi _5532__128 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net128));
 sg13g2_tiehi _5284__129 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net129));
 sg13g2_tiehi _5440__130 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net130));
 sg13g2_tiehi _5283__131 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net131));
 sg13g2_tiehi _5282__132 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net132));
 sg13g2_tiehi _5562__133 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net133));
 sg13g2_tiehi _5281__134 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net134));
 sg13g2_tiehi _5439__135 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net135));
 sg13g2_tiehi _5280__136 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net136));
 sg13g2_tiehi _5531__137 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net137));
 sg13g2_tiehi _5279__138 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net138));
 sg13g2_tiehi _5438__139 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net139));
 sg13g2_tiehi _5278__140 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net140));
 sg13g2_tiehi _5561__141 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net141));
 sg13g2_tiehi _5277__142 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net142));
 sg13g2_tiehi _5437__143 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net143));
 sg13g2_tiehi _5276__144 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net144));
 sg13g2_tiehi _5530__145 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net145));
 sg13g2_tiehi _5275__146 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net146));
 sg13g2_tiehi _5436__147 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net147));
 sg13g2_tiehi _5274__148 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net148));
 sg13g2_tiehi _5560__149 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net149));
 sg13g2_tiehi _5273__150 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net150));
 sg13g2_tiehi _5435__151 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net151));
 sg13g2_tiehi _5272__152 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net152));
 sg13g2_tiehi _5529__153 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net153));
 sg13g2_tiehi _5271__154 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net154));
 sg13g2_tiehi _5434__155 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net155));
 sg13g2_tiehi _5270__156 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net156));
 sg13g2_tiehi _5559__157 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net157));
 sg13g2_tiehi _5269__158 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net158));
 sg13g2_tiehi _5433__159 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net159));
 sg13g2_tiehi _5268__160 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net160));
 sg13g2_tiehi _5528__161 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net161));
 sg13g2_tiehi _5267__162 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net162));
 sg13g2_tiehi _5432__163 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net163));
 sg13g2_tiehi _5266__164 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net164));
 sg13g2_tiehi _5527__165 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net165));
 sg13g2_tiehi _5265__166 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net166));
 sg13g2_tiehi _5431__167 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net167));
 sg13g2_tiehi _5264__168 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net168));
 sg13g2_tiehi _5526__169 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net169));
 sg13g2_tiehi _5263__170 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net170));
 sg13g2_tiehi _5430__171 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net171));
 sg13g2_tiehi _5262__172 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net172));
 sg13g2_tiehi _5261__173 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net173));
 sg13g2_tiehi _5525__174 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net174));
 sg13g2_tiehi _5260__175 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net175));
 sg13g2_tiehi _5429__176 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net176));
 sg13g2_tiehi _5259__177 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net177));
 sg13g2_tiehi _5524__178 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net178));
 sg13g2_tiehi _5258__179 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net179));
 sg13g2_tiehi _5428__180 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net180));
 sg13g2_tiehi _5257__181 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net181));
 sg13g2_tiehi _5523__182 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net182));
 sg13g2_tiehi _5256__183 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net183));
 sg13g2_tiehi _5427__184 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net184));
 sg13g2_tiehi _5255__185 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net185));
 sg13g2_tiehi _5522__186 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net186));
 sg13g2_tiehi _5254__187 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net187));
 sg13g2_tiehi _5426__188 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net188));
 sg13g2_tiehi _5253__189 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net189));
 sg13g2_tiehi _5521__190 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net190));
 sg13g2_tiehi _5252__191 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net191));
 sg13g2_tiehi _5425__192 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net192));
 sg13g2_tiehi _5251__193 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net193));
 sg13g2_tiehi _5558__194 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net194));
 sg13g2_tiehi _5250__195 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net195));
 sg13g2_tiehi _5424__196 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net196));
 sg13g2_tiehi _5249__197 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net197));
 sg13g2_tiehi _5520__198 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net198));
 sg13g2_tiehi _5248__199 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net199));
 sg13g2_tiehi _5423__200 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net200));
 sg13g2_tiehi _5247__201 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net201));
 sg13g2_tiehi _5557__202 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net202));
 sg13g2_tiehi _5246__203 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net203));
 sg13g2_tiehi _5422__204 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net204));
 sg13g2_tiehi _5245__205 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net205));
 sg13g2_tiehi _5519__206 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net206));
 sg13g2_tiehi _5244__207 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net207));
 sg13g2_tiehi _5421__208 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net208));
 sg13g2_tiehi _5243__209 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net209));
 sg13g2_tiehi _5556__210 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net210));
 sg13g2_tiehi _5242__211 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net211));
 sg13g2_tiehi _5420__212 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net212));
 sg13g2_tiehi _5518__213 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net213));
 sg13g2_tiehi _5419__214 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net214));
 sg13g2_tiehi _5555__215 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net215));
 sg13g2_tiehi _5418__216 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net216));
 sg13g2_tiehi _5517__217 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net217));
 sg13g2_tiehi _5417__218 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net218));
 sg13g2_tiehi _5554__219 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net219));
 sg13g2_tiehi _5416__220 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net220));
 sg13g2_tiehi _5516__221 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net221));
 sg13g2_tiehi _5415__222 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net222));
 sg13g2_tiehi _5305__223 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net223));
 sg13g2_tiehi _5414__224 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net224));
 sg13g2_tiehi _5515__225 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net225));
 sg13g2_tiehi _5413__226 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net226));
 sg13g2_tiehi _5553__227 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net227));
 sg13g2_tiehi _5412__228 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net228));
 sg13g2_tiehi _5514__229 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net229));
 sg13g2_tiehi _5411__230 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net230));
 sg13g2_tiehi _5583__231 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net231));
 sg13g2_tiehi _5410__232 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net232));
 sg13g2_tiehi _5513__233 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net233));
 sg13g2_tiehi _5409__234 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net234));
 sg13g2_tiehi _5552__235 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net235));
 sg13g2_tiehi _5408__236 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net236));
 sg13g2_tiehi _5512__237 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net237));
 sg13g2_tiehi _5407__238 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net238));
 sg13g2_tiehi _5582__239 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net239));
 sg13g2_tiehi _5406__240 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net240));
 sg13g2_tiehi _5511__241 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net241));
 sg13g2_tiehi _5405__242 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net242));
 sg13g2_tiehi _5551__243 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net243));
 sg13g2_tiehi _5404__244 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net244));
 sg13g2_tiehi _5510__245 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net245));
 sg13g2_tiehi _5403__246 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net246));
 sg13g2_tiehi _5581__247 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net247));
 sg13g2_tiehi _5402__248 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net248));
 sg13g2_tiehi _5509__249 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net249));
 sg13g2_tiehi _5401__250 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net250));
 sg13g2_tiehi _5550__251 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net251));
 sg13g2_tiehi _5400__252 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net252));
 sg13g2_tiehi _5508__253 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net253));
 sg13g2_tiehi _5399__254 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net254));
 sg13g2_tiehi _5580__255 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net255));
 sg13g2_tiehi _5398__256 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net256));
 sg13g2_tiehi _5507__257 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net257));
 sg13g2_tiehi _5397__258 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net258));
 sg13g2_tiehi _5549__259 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net259));
 sg13g2_tiehi _5396__260 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net260));
 sg13g2_tiehi _5506__261 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net261));
 sg13g2_tiehi _5395__262 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net262));
 sg13g2_tiehi _5579__263 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net263));
 sg13g2_tiehi _5394__264 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net264));
 sg13g2_tiehi _5505__265 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net265));
 sg13g2_tiehi _5393__266 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net266));
 sg13g2_tiehi _5504__267 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net267));
 sg13g2_tiehi _5392__268 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net268));
 sg13g2_tiehi _5503__269 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net269));
 sg13g2_tiehi _5391__270 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net270));
 sg13g2_tiehi _5502__271 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net271));
 sg13g2_tiehi _5390__272 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net272));
 sg13g2_tiehi _5501__273 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net273));
 sg13g2_tiehi _5389__274 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net274));
 sg13g2_tiehi _5500__275 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net275));
 sg13g2_tiehi _5388__276 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net276));
 sg13g2_tiehi _5499__277 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net277));
 sg13g2_tiehi _5387__278 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net278));
 sg13g2_tiehi _5498__279 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net279));
 sg13g2_tiehi _5386__280 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net280));
 sg13g2_tiehi _5497__281 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net281));
 sg13g2_tiehi _5385__282 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net282));
 sg13g2_tiehi _5496__283 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net283));
 sg13g2_tiehi _5384__284 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net284));
 sg13g2_tiehi _5548__285 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net285));
 sg13g2_tiehi _5383__286 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net286));
 sg13g2_tiehi _5495__287 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net287));
 sg13g2_tiehi _5382__288 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net288));
 sg13g2_tiehi _5578__289 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net289));
 sg13g2_tiehi _5381__290 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net290));
 sg13g2_tiehi _5494__291 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net291));
 sg13g2_tiehi _5380__292 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net292));
 sg13g2_tiehi _5547__293 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net293));
 sg13g2_tiehi _5379__294 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net294));
 sg13g2_tiehi _5493__295 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net295));
 sg13g2_tiehi _5378__296 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net296));
 sg13g2_tiehi _5492__297 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net297));
 sg13g2_tiehi _5377__298 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net298));
 sg13g2_tiehi _5491__299 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net299));
 sg13g2_tiehi _5376__300 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net300));
 sg13g2_tiehi _5490__301 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net301));
 sg13g2_tiehi _5375__302 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net302));
 sg13g2_tiehi _5489__303 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net303));
 sg13g2_tiehi _5374__304 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net304));
 sg13g2_tiehi _5488__305 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net305));
 sg13g2_tiehi _5373__306 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net306));
 sg13g2_tiehi _5577__307 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net307));
 sg13g2_tiehi _5372__308 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net308));
 sg13g2_tiehi _5487__309 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net309));
 sg13g2_tiehi _5371__310 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net310));
 sg13g2_tiehi _5486__311 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net311));
 sg13g2_tiehi _5370__312 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net312));
 sg13g2_tiehi _5546__313 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net313));
 sg13g2_tiehi _5369__314 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net314));
 sg13g2_tiehi _5485__315 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net315));
 sg13g2_tiehi _5368__316 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net316));
 sg13g2_tiehi _5484__317 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net317));
 sg13g2_tiehi _5367__318 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net318));
 sg13g2_tiehi _5483__319 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net319));
 sg13g2_tiehi _5366__320 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net320));
 sg13g2_tiehi _5482__321 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net321));
 sg13g2_tiehi _5365__322 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net322));
 sg13g2_tiehi _5481__323 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net323));
 sg13g2_tiehi _5364__324 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net324));
 sg13g2_tiehi _5480__325 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net325));
 sg13g2_tiehi _5363__326 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net326));
 sg13g2_tiehi _5479__327 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net327));
 sg13g2_tiehi _5362__328 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net328));
 sg13g2_tiehi _5478__329 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net329));
 sg13g2_tiehi _5361__330 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net330));
 sg13g2_tiehi _5477__331 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net331));
 sg13g2_tiehi _5360__332 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net332));
 sg13g2_tiehi _5476__333 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net333));
 sg13g2_tiehi _5359__334 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net334));
 sg13g2_tiehi _5475__335 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net335));
 sg13g2_tiehi _5358__336 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net336));
 sg13g2_tiehi _5474__337 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net337));
 sg13g2_tiehi _5357__338 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net338));
 sg13g2_tiehi _5473__339 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net339));
 sg13g2_tiehi _5356__340 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net340));
 sg13g2_tiehi _5472__341 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net341));
 sg13g2_tiehi _5355__342 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net342));
 sg13g2_tiehi _5471__343 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net343));
 sg13g2_tiehi _5354__344 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net344));
 sg13g2_tiehi _5470__345 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net345));
 sg13g2_tiehi _5353__346 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net346));
 sg13g2_tiehi _5469__347 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net347));
 sg13g2_tiehi _5352__348 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net348));
 sg13g2_tiehi _5468__349 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net349));
 sg13g2_tiehi _5351__350 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net350));
 sg13g2_tiehi _5576__351 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net351));
 sg13g2_tiehi _5350__352 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net352));
 sg13g2_tiehi _5467__353 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net353));
 sg13g2_tiehi _5349__354 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net354));
 sg13g2_tiehi _5545__355 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net355));
 sg13g2_tiehi _5348__356 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net356));
 sg13g2_tiehi _5466__357 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net357));
 sg13g2_tiehi _5347__358 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net358));
 sg13g2_tiehi _5575__359 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net359));
 sg13g2_tiehi _5346__360 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net360));
 sg13g2_tiehi _5465__361 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net361));
 sg13g2_tiehi _5345__362 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net362));
 sg13g2_tiehi _5544__363 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net363));
 sg13g2_tiehi _5344__364 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net364));
 sg13g2_tiehi _5464__365 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net365));
 sg13g2_tiehi _5343__366 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net366));
 sg13g2_tiehi _5574__367 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net367));
 sg13g2_tiehi _5342__368 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net368));
 sg13g2_tiehi _5463__369 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net369));
 sg13g2_tiehi _5341__370 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net370));
 sg13g2_tiehi _5340__371 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net371));
 sg13g2_tiehi _5339__372 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net372));
 sg13g2_buf_8 clkbuf_leaf_0_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_tiny_wrapper_9 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net9));
 sg13g2_tielo heichips25_tiny_wrapper_10 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net10));
 sg13g2_tielo heichips25_tiny_wrapper_11 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net11));
 sg13g2_tielo heichips25_tiny_wrapper_12 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net12));
 sg13g2_tielo heichips25_tiny_wrapper_13 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net13));
 sg13g2_tielo heichips25_tiny_wrapper_14 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net14));
 sg13g2_tielo heichips25_tiny_wrapper_15 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net15));
 sg13g2_tielo heichips25_tiny_wrapper_16 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net16));
 sg13g2_tielo heichips25_tiny_wrapper_17 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net17));
 sg13g2_tielo heichips25_tiny_wrapper_18 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net18));
 sg13g2_tielo heichips25_tiny_wrapper_19 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net19));
 sg13g2_tielo heichips25_tiny_wrapper_20 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net20));
 sg13g2_tielo heichips25_tiny_wrapper_21 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net21));
 sg13g2_tielo heichips25_tiny_wrapper_22 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net22));
 sg13g2_tielo heichips25_tiny_wrapper_23 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net23));
 sg13g2_tielo heichips25_tiny_wrapper_24 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net24));
 sg13g2_tielo heichips25_tiny_wrapper_25 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net25));
 sg13g2_tielo heichips25_tiny_wrapper_26 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net26));
 sg13g2_tielo heichips25_tiny_wrapper_27 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net27));
 sg13g2_tielo heichips25_tiny_wrapper_28 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net28));
 sg13g2_tielo heichips25_tiny_wrapper_29 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net29));
 sg13g2_tiehi _5338__30 (.VDD(VPWR),
    .VSS(VGND),
    .L_HI(net30));
 sg13g2_buf_2 _5949_ (.A(\falu_i.falutop.i2c_inst.sda_o ),
    .X(net6),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 _5950_ (.A(\ppwm_i.u_ppwm.data_o ),
    .X(net7),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout563 (.A(net564),
    .X(net563),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout564 (.A(net565),
    .X(net564),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout565 (.A(_1278_),
    .X(net565),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout566 (.A(_1278_),
    .X(net566),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout567 (.A(net568),
    .X(net567),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout568 (.A(_1132_),
    .X(net568),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout569 (.A(_0814_),
    .X(net569),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout570 (.A(_0814_),
    .X(net570),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout571 (.A(_0628_),
    .X(net571),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout572 (.A(net573),
    .X(net572),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout573 (.A(_0615_),
    .X(net573),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout574 (.A(_0649_),
    .X(net574),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout575 (.A(_0617_),
    .X(net575),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout576 (.A(_0617_),
    .X(net576),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout577 (.A(net580),
    .X(net577),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout578 (.A(net580),
    .X(net578),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout579 (.A(net580),
    .X(net579),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout580 (.A(_0608_),
    .X(net580),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout581 (.A(net583),
    .X(net581),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout582 (.A(net583),
    .X(net582),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout583 (.A(_0530_),
    .X(net583),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout584 (.A(net585),
    .X(net584),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout585 (.A(_2390_),
    .X(net585),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout586 (.A(_2375_),
    .X(net586),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout587 (.A(_1295_),
    .X(net587),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout588 (.A(net590),
    .X(net588),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout589 (.A(net590),
    .X(net589),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout590 (.A(_0610_),
    .X(net590),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout591 (.A(net592),
    .X(net591),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout592 (.A(net593),
    .X(net592),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout593 (.A(net597),
    .X(net593),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout594 (.A(net596),
    .X(net594),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout595 (.A(net596),
    .X(net595),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout596 (.A(net597),
    .X(net596),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout597 (.A(_2404_),
    .X(net597),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout598 (.A(net599),
    .X(net598),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout599 (.A(_2404_),
    .X(net599),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout600 (.A(net604),
    .X(net600),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout601 (.A(net604),
    .X(net601),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout602 (.A(net604),
    .X(net602),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout603 (.A(net604),
    .X(net603),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout604 (.A(_2374_),
    .X(net604),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout605 (.A(net606),
    .X(net605),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout606 (.A(_1106_),
    .X(net606),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout607 (.A(_1105_),
    .X(net607),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout608 (.A(_2418_),
    .X(net608),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout609 (.A(net610),
    .X(net609),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout610 (.A(_2389_),
    .X(net610),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout611 (.A(net613),
    .X(net611),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout612 (.A(net613),
    .X(net612),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout613 (.A(_2389_),
    .X(net613),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout614 (.A(_1590_),
    .X(net614),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout615 (.A(_1317_),
    .X(net615),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout616 (.A(_1281_),
    .X(net616),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout617 (.A(net621),
    .X(net617),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout618 (.A(net621),
    .X(net618),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout619 (.A(net621),
    .X(net619),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout620 (.A(net621),
    .X(net620),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout621 (.A(_1136_),
    .X(net621),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout622 (.A(_1078_),
    .X(net622),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout623 (.A(net624),
    .X(net623),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout624 (.A(net626),
    .X(net624),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout625 (.A(net626),
    .X(net625),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout626 (.A(_1077_),
    .X(net626),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout627 (.A(net629),
    .X(net627),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout628 (.A(net629),
    .X(net628),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout629 (.A(_1076_),
    .X(net629),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout630 (.A(_1075_),
    .X(net630),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout631 (.A(_1306_),
    .X(net631),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout632 (.A(_1242_),
    .X(net632),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout633 (.A(net635),
    .X(net633),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout634 (.A(net635),
    .X(net634),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout635 (.A(_1134_),
    .X(net635),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout636 (.A(net637),
    .X(net636),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout637 (.A(_1134_),
    .X(net637),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout638 (.A(net640),
    .X(net638),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout639 (.A(net640),
    .X(net639),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout640 (.A(_1073_),
    .X(net640),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout641 (.A(net642),
    .X(net641),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout642 (.A(net645),
    .X(net642),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout643 (.A(net645),
    .X(net643),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout644 (.A(net645),
    .X(net644),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout645 (.A(net651),
    .X(net645),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout646 (.A(net651),
    .X(net646),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout647 (.A(net651),
    .X(net647),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout648 (.A(net650),
    .X(net648),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout649 (.A(net650),
    .X(net649),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout650 (.A(net651),
    .X(net650),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout651 (.A(net652),
    .X(net651),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout652 (.A(_0908_),
    .X(net652),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout653 (.A(net655),
    .X(net653),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout654 (.A(net655),
    .X(net654),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout655 (.A(net666),
    .X(net655),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout656 (.A(net658),
    .X(net656),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout657 (.A(net658),
    .X(net657),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout658 (.A(net666),
    .X(net658),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout659 (.A(net663),
    .X(net659),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout660 (.A(net663),
    .X(net660),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout661 (.A(net663),
    .X(net661),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout662 (.A(net663),
    .X(net662),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout663 (.A(net666),
    .X(net663),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout664 (.A(net665),
    .X(net664),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout665 (.A(net666),
    .X(net665),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout666 (.A(net680),
    .X(net666),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout667 (.A(net668),
    .X(net667),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout668 (.A(net679),
    .X(net668),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout669 (.A(net670),
    .X(net669),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout670 (.A(net671),
    .X(net670),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout671 (.A(net679),
    .X(net671),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout672 (.A(net675),
    .X(net672),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout673 (.A(net675),
    .X(net673),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout674 (.A(net675),
    .X(net674),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout675 (.A(net679),
    .X(net675),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout676 (.A(net678),
    .X(net676),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout677 (.A(net678),
    .X(net677),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout678 (.A(net679),
    .X(net678),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout679 (.A(net680),
    .X(net679),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout680 (.A(net884),
    .X(net680),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout681 (.A(net683),
    .X(net681),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout682 (.A(net683),
    .X(net682),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout683 (.A(_0386_),
    .X(net683),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout684 (.A(net687),
    .X(net684),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout685 (.A(net687),
    .X(net685),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout686 (.A(net687),
    .X(net686),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout687 (.A(_0902_),
    .X(net687),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout688 (.A(_2312_),
    .X(net688),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout689 (.A(_2312_),
    .X(net689),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout690 (.A(net691),
    .X(net690),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout691 (.A(_2312_),
    .X(net691),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout692 (.A(_2311_),
    .X(net692),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout693 (.A(_2311_),
    .X(net693),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout694 (.A(net695),
    .X(net694),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout695 (.A(_2311_),
    .X(net695),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout696 (.A(net699),
    .X(net696),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout697 (.A(net698),
    .X(net697),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout698 (.A(net699),
    .X(net698),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout699 (.A(_2309_),
    .X(net699),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout700 (.A(net701),
    .X(net700),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout701 (.A(net704),
    .X(net701),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout702 (.A(net703),
    .X(net702),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout703 (.A(net704),
    .X(net703),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout704 (.A(_2306_),
    .X(net704),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout705 (.A(_2302_),
    .X(net705),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout706 (.A(_2302_),
    .X(net706),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout707 (.A(_2295_),
    .X(net707),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout708 (.A(_2256_),
    .X(net708),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout709 (.A(_2256_),
    .X(net709),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout710 (.A(net715),
    .X(net710),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout711 (.A(net713),
    .X(net711),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout712 (.A(net713),
    .X(net712),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout713 (.A(net714),
    .X(net713),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout714 (.A(net715),
    .X(net714),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout715 (.A(\falu_i.falutop.alu_data_in[15] ),
    .X(net715),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout716 (.A(net717),
    .X(net716),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout717 (.A(net720),
    .X(net717),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout718 (.A(net719),
    .X(net718),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout719 (.A(net720),
    .X(net719),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout720 (.A(\falu_i.falutop.alu_data_in[14] ),
    .X(net720),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout721 (.A(net722),
    .X(net721),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout722 (.A(\falu_i.falutop.alu_data_in[13] ),
    .X(net722),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout723 (.A(net724),
    .X(net723),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout724 (.A(\falu_i.falutop.alu_data_in[13] ),
    .X(net724),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout725 (.A(net726),
    .X(net725),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout726 (.A(\falu_i.falutop.alu_data_in[12] ),
    .X(net726),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout727 (.A(net729),
    .X(net727),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout728 (.A(net729),
    .X(net728),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout729 (.A(\falu_i.falutop.alu_data_in[12] ),
    .X(net729),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout730 (.A(\falu_i.falutop.alu_data_in[11] ),
    .X(net730),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout731 (.A(\falu_i.falutop.alu_data_in[11] ),
    .X(net731),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout732 (.A(net733),
    .X(net732),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout733 (.A(net734),
    .X(net733),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout734 (.A(\falu_i.falutop.alu_data_in[11] ),
    .X(net734),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout735 (.A(net736),
    .X(net735),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout736 (.A(net739),
    .X(net736),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout737 (.A(net738),
    .X(net737),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout738 (.A(net739),
    .X(net738),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout739 (.A(\falu_i.falutop.alu_data_in[10] ),
    .X(net739),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout740 (.A(\falu_i.falutop.alu_data_in[9] ),
    .X(net740),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout741 (.A(net742),
    .X(net741),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout742 (.A(\falu_i.falutop.alu_data_in[9] ),
    .X(net742),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout743 (.A(net746),
    .X(net743),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout744 (.A(net746),
    .X(net744),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout745 (.A(net746),
    .X(net745),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout746 (.A(\falu_i.falutop.alu_data_in[8] ),
    .X(net746),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout747 (.A(net748),
    .X(net747),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout748 (.A(net749),
    .X(net748),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout749 (.A(net1131),
    .X(net749),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout750 (.A(\falu_i.falutop.alu_data_in[5] ),
    .X(net750),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout751 (.A(\falu_i.falutop.alu_data_in[5] ),
    .X(net751),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout752 (.A(net754),
    .X(net752),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout753 (.A(net754),
    .X(net753),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout754 (.A(\falu_i.falutop.alu_data_in[4] ),
    .X(net754),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout755 (.A(net758),
    .X(net755),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout756 (.A(net757),
    .X(net756),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout757 (.A(net758),
    .X(net757),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout758 (.A(net759),
    .X(net758),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout759 (.A(net760),
    .X(net759),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout760 (.A(\falu_i.falutop.alu_data_in[3] ),
    .X(net760),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout761 (.A(net764),
    .X(net761),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout762 (.A(net763),
    .X(net762),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout763 (.A(net764),
    .X(net763),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout764 (.A(net765),
    .X(net764),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout765 (.A(\falu_i.falutop.alu_data_in[2] ),
    .X(net765),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout766 (.A(net767),
    .X(net766),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout767 (.A(\falu_i.falutop.alu_data_in[1] ),
    .X(net767),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout768 (.A(net769),
    .X(net768),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout769 (.A(net770),
    .X(net769),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout770 (.A(\falu_i.falutop.alu_data_in[0] ),
    .X(net770),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout771 (.A(net964),
    .X(net771),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout772 (.A(net938),
    .X(net772),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout773 (.A(net774),
    .X(net773),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout774 (.A(net775),
    .X(net774),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout775 (.A(net776),
    .X(net775),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout776 (.A(net1178),
    .X(net776),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout777 (.A(\falu_i.falutop.data_in[7] ),
    .X(net777),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout778 (.A(net779),
    .X(net778),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout779 (.A(net887),
    .X(net779),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout780 (.A(net887),
    .X(net780),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout781 (.A(\falu_i.falutop.div_inst.start ),
    .X(net781),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout782 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .X(net782),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout783 (.A(net1194),
    .X(net783),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout784 (.A(net785),
    .X(net784),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout785 (.A(net1196),
    .X(net785),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout786 (.A(net1192),
    .X(net786),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout787 (.A(\ppwm_i.u_ppwm.pc[3] ),
    .X(net787),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout788 (.A(net790),
    .X(net788),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout789 (.A(net790),
    .X(net789),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout790 (.A(net1193),
    .X(net790),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout791 (.A(net1168),
    .X(net791),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout792 (.A(\ppwm_i.u_ppwm.pc[1] ),
    .X(net792),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout793 (.A(\ppwm_i.u_ppwm.pc[0] ),
    .X(net793),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout794 (.A(\ppwm_i.u_ppwm.pc[0] ),
    .X(net794),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout795 (.A(net796),
    .X(net795),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout796 (.A(net797),
    .X(net796),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout797 (.A(_2294_),
    .X(net797),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout798 (.A(net799),
    .X(net798),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout799 (.A(_2294_),
    .X(net799),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout800 (.A(_2289_),
    .X(net800),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout801 (.A(_2289_),
    .X(net801),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout802 (.A(_2289_),
    .X(net802),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout803 (.A(net805),
    .X(net803),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout804 (.A(net805),
    .X(net804),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout805 (.A(net806),
    .X(net805),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout806 (.A(net814),
    .X(net806),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout807 (.A(net808),
    .X(net807),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout808 (.A(net811),
    .X(net808),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout809 (.A(net811),
    .X(net809),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout810 (.A(net811),
    .X(net810),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout811 (.A(net814),
    .X(net811),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout812 (.A(net814),
    .X(net812),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout813 (.A(net814),
    .X(net813),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout814 (.A(rst_n),
    .X(net814),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout815 (.A(net817),
    .X(net815),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout816 (.A(net817),
    .X(net816),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout817 (.A(net823),
    .X(net817),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout818 (.A(net820),
    .X(net818),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout819 (.A(net820),
    .X(net819),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout820 (.A(net823),
    .X(net820),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout821 (.A(net822),
    .X(net821),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout822 (.A(net823),
    .X(net822),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout823 (.A(rst_n),
    .X(net823),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout824 (.A(net832),
    .X(net824),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout825 (.A(net826),
    .X(net825),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout826 (.A(net832),
    .X(net826),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout827 (.A(net831),
    .X(net827),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout828 (.A(net831),
    .X(net828),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout829 (.A(net830),
    .X(net829),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout830 (.A(net831),
    .X(net830),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout831 (.A(net832),
    .X(net831),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_2 fanout832 (.A(net833),
    .X(net832),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 fanout833 (.A(net842),
    .X(net833),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout834 (.A(net835),
    .X(net834),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout835 (.A(net842),
    .X(net835),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout836 (.A(net842),
    .X(net836),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout837 (.A(net838),
    .X(net837),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout838 (.A(net841),
    .X(net838),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout839 (.A(net840),
    .X(net839),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout840 (.A(net841),
    .X(net840),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout841 (.A(net842),
    .X(net841),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 fanout842 (.A(rst_n),
    .X(net842),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input3 (.A(ui_in[3]),
    .X(net3),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input4 (.A(ui_in[4]),
    .X(net4),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 input5 (.A(ui_in[5]),
    .X(net5),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output6 (.A(net6),
    .X(uo_out[0]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_1 output7 (.A(net7),
    .X(uo_out[4]),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_tielo heichips25_tiny_wrapper_8 (.VDD(VPWR),
    .VSS(VGND),
    .L_LO(net8));
 sg13g2_buf_8 clkbuf_leaf_1_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_1_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_2_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_2_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_3_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_3_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_4_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_4_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_5_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_5_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_6_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_6_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_7_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_7_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_8_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_8_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_9_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_9_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_10_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_10_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_11_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_11_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_12_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_12_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_13_clk (.A(clknet_3_3__leaf_clk),
    .X(clknet_leaf_13_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_14_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_14_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_15_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_15_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_16_clk (.A(clknet_3_2__leaf_clk),
    .X(clknet_leaf_16_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_17_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_17_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_18_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_19_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_19_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_20_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_20_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_21_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_21_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_22_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_22_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_23_clk (.A(clknet_3_4__leaf_clk),
    .X(clknet_leaf_23_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_24_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_24_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_25_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_25_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_26_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_26_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_27_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_27_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_28_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_28_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_29_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_29_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_30_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_30_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_31_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_31_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_32_clk (.A(clknet_3_7__leaf_clk),
    .X(clknet_leaf_32_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_33_clk (.A(clknet_3_6__leaf_clk),
    .X(clknet_leaf_33_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_34_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_34_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_35_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_36_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_37_clk (.A(clknet_3_5__leaf_clk),
    .X(clknet_leaf_37_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_38_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_38_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_39_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_39_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_40_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_40_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_41_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_41_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_42_clk (.A(clknet_3_1__leaf_clk),
    .X(clknet_leaf_42_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_43_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_43_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_leaf_44_clk (.A(clknet_3_0__leaf_clk),
    .X(clknet_leaf_44_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_0__f_clk (.A(clknet_0_clk),
    .X(clknet_3_0__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_1__f_clk (.A(clknet_0_clk),
    .X(clknet_3_1__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_2__f_clk (.A(clknet_0_clk),
    .X(clknet_3_2__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_3__f_clk (.A(clknet_0_clk),
    .X(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_4__f_clk (.A(clknet_0_clk),
    .X(clknet_3_4__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_5__f_clk (.A(clknet_0_clk),
    .X(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_6__f_clk (.A(clknet_0_clk),
    .X(clknet_3_6__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkbuf_3_7__f_clk (.A(clknet_0_clk),
    .X(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload0 (.A(clknet_3_3__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload1 (.A(clknet_3_5__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_buf_8 clkload2 (.A(clknet_3_7__leaf_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_1 clkload3 (.VDD(VPWR),
    .A(clknet_leaf_44_clk),
    .VSS(VGND));
 sg13g2_inv_8 clkload4 (.A(clknet_leaf_18_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_4 clkload5 (.A(clknet_leaf_35_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_inv_8 clkload6 (.A(clknet_leaf_36_clk),
    .VDD(VPWR),
    .VSS(VGND));
 sg13g2_dlygate4sd3_1 hold1 (.A(\ppwm_i.u_ppwm.u_mem.data_sync1 ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net373));
 sg13g2_dlygate4sd3_1 hold2 (.A(\ppwm_i.u_ppwm.u_mem.clk_prog_sync1 ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net374));
 sg13g2_dlygate4sd3_1 hold3 (.A(\ppwm_i.u_ppwm.u_mem.clk_prog_sync2 ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net375));
 sg13g2_dlygate4sd3_1 hold4 (.A(\ppwm_i.u_ppwm.polarity ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net376));
 sg13g2_dlygate4sd3_1 hold5 (.A(_0065_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net377));
 sg13g2_dlygate4sd3_1 hold6 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net378));
 sg13g2_dlygate4sd3_1 hold7 (.A(_0212_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net379));
 sg13g2_dlygate4sd3_1 hold8 (.A(\falu_i.falutop.div_inst.done ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net380));
 sg13g2_dlygate4sd3_1 hold9 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net381));
 sg13g2_dlygate4sd3_1 hold10 (.A(_0024_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net382));
 sg13g2_dlygate4sd3_1 hold11 (.A(\ppwm_i.u_ppwm.u_mem.memory[75] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net383));
 sg13g2_dlygate4sd3_1 hold12 (.A(_0174_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net384));
 sg13g2_dlygate4sd3_1 hold13 (.A(\ppwm_i.u_ppwm.u_ex.state_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net385));
 sg13g2_dlygate4sd3_1 hold14 (.A(_2426_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net386));
 sg13g2_dlygate4sd3_1 hold15 (.A(_0001_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net387));
 sg13g2_dlygate4sd3_1 hold16 (.A(\falu_i.falutop.div_inst.a[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net388));
 sg13g2_dlygate4sd3_1 hold17 (.A(_0337_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net389));
 sg13g2_dlygate4sd3_1 hold18 (.A(\ppwm_i.u_ppwm.u_mem.memory[92] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net390));
 sg13g2_dlygate4sd3_1 hold19 (.A(_0191_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net391));
 sg13g2_dlygate4sd3_1 hold20 (.A(\ppwm_i.u_ppwm.u_mem.memory[103] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net392));
 sg13g2_dlygate4sd3_1 hold21 (.A(_0202_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net393));
 sg13g2_dlygate4sd3_1 hold22 (.A(\ppwm_i.u_ppwm.u_mem.memory[56] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net394));
 sg13g2_dlygate4sd3_1 hold23 (.A(_0156_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net395));
 sg13g2_dlygate4sd3_1 hold24 (.A(\falu_i.falutop.div_inst.acc_next[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net396));
 sg13g2_dlygate4sd3_1 hold25 (.A(_0286_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net397));
 sg13g2_dlygate4sd3_1 hold26 (.A(\ppwm_i.u_ppwm.u_mem.memory[55] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net398));
 sg13g2_dlygate4sd3_1 hold27 (.A(\falu_i.falutop.div_inst.quo[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net399));
 sg13g2_dlygate4sd3_1 hold28 (.A(_0280_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net400));
 sg13g2_dlygate4sd3_1 hold29 (.A(\ppwm_i.u_ppwm.u_mem.memory[93] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net401));
 sg13g2_dlygate4sd3_1 hold30 (.A(\ppwm_i.u_ppwm.u_mem.memory[24] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net402));
 sg13g2_dlygate4sd3_1 hold31 (.A(_0123_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net403));
 sg13g2_dlygate4sd3_1 hold32 (.A(\ppwm_i.u_ppwm.u_mem.memory[76] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net404));
 sg13g2_dlygate4sd3_1 hold33 (.A(\falu_i.falutop.div_inst.quo[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net405));
 sg13g2_dlygate4sd3_1 hold34 (.A(_0283_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net406));
 sg13g2_dlygate4sd3_1 hold35 (.A(\ppwm_i.u_ppwm.u_mem.memory[50] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net407));
 sg13g2_dlygate4sd3_1 hold36 (.A(_0150_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net408));
 sg13g2_dlygate4sd3_1 hold37 (.A(\falu_i.falutop.div_inst.i[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net409));
 sg13g2_dlygate4sd3_1 hold38 (.A(_0254_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net410));
 sg13g2_dlygate4sd3_1 hold39 (.A(\falu_i.falutop.div_inst.quo[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net411));
 sg13g2_dlygate4sd3_1 hold40 (.A(_0281_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net412));
 sg13g2_dlygate4sd3_1 hold41 (.A(\falu_i.falutop.div_inst.b[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net413));
 sg13g2_dlygate4sd3_1 hold42 (.A(_0330_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net414));
 sg13g2_dlygate4sd3_1 hold43 (.A(\ppwm_i.u_ppwm.u_mem.memory[71] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net415));
 sg13g2_dlygate4sd3_1 hold44 (.A(_0170_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net416));
 sg13g2_dlygate4sd3_1 hold45 (.A(\ppwm_i.u_ppwm.u_mem.memory[82] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net417));
 sg13g2_dlygate4sd3_1 hold46 (.A(_0181_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net418));
 sg13g2_dlygate4sd3_1 hold47 (.A(\ppwm_i.u_ppwm.u_ex.state_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net419));
 sg13g2_dlygate4sd3_1 hold48 (.A(\falu_i.falutop.i2c_inst.op[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net420));
 sg13g2_dlygate4sd3_1 hold49 (.A(_0092_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net421));
 sg13g2_dlygate4sd3_1 hold50 (.A(\ppwm_i.u_ppwm.u_mem.memory[39] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net422));
 sg13g2_dlygate4sd3_1 hold51 (.A(_0138_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net423));
 sg13g2_dlygate4sd3_1 hold52 (.A(\ppwm_i.u_ppwm.u_mem.memory[37] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net424));
 sg13g2_dlygate4sd3_1 hold53 (.A(_0137_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net425));
 sg13g2_dlygate4sd3_1 hold54 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net426));
 sg13g2_dlygate4sd3_1 hold55 (.A(_0029_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net427));
 sg13g2_dlygate4sd3_1 hold56 (.A(\falu_i.falutop.i2c_inst.op[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net428));
 sg13g2_dlygate4sd3_1 hold57 (.A(_0095_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net429));
 sg13g2_dlygate4sd3_1 hold58 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net430));
 sg13g2_dlygate4sd3_1 hold59 (.A(_0031_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net431));
 sg13g2_dlygate4sd3_1 hold60 (.A(\falu_i.falutop.div_inst.quo[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net432));
 sg13g2_dlygate4sd3_1 hold61 (.A(_0284_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net433));
 sg13g2_dlygate4sd3_1 hold62 (.A(\ppwm_i.u_ppwm.u_mem.memory[49] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net434));
 sg13g2_dlygate4sd3_1 hold63 (.A(\falu_i.falutop.div_inst.quo[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net435));
 sg13g2_dlygate4sd3_1 hold64 (.A(_0282_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net436));
 sg13g2_dlygate4sd3_1 hold65 (.A(\ppwm_i.u_ppwm.u_mem.memory[61] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net437));
 sg13g2_dlygate4sd3_1 hold66 (.A(_0160_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net438));
 sg13g2_dlygate4sd3_1 hold67 (.A(\falu_i.falutop.div_inst.a[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net439));
 sg13g2_dlygate4sd3_1 hold68 (.A(_0342_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net440));
 sg13g2_dlygate4sd3_1 hold69 (.A(\ppwm_i.u_ppwm.u_mem.memory[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net441));
 sg13g2_dlygate4sd3_1 hold70 (.A(_0108_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net442));
 sg13g2_dlygate4sd3_1 hold71 (.A(\ppwm_i.u_ppwm.u_mem.memory[53] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net443));
 sg13g2_dlygate4sd3_1 hold72 (.A(_0152_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net444));
 sg13g2_dlygate4sd3_1 hold73 (.A(\ppwm_i.u_ppwm.u_mem.memory[107] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net445));
 sg13g2_dlygate4sd3_1 hold74 (.A(_0206_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net446));
 sg13g2_dlygate4sd3_1 hold75 (.A(\ppwm_i.u_ppwm.u_mem.memory[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net447));
 sg13g2_dlygate4sd3_1 hold76 (.A(_0116_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net448));
 sg13g2_dlygate4sd3_1 hold77 (.A(\ppwm_i.u_ppwm.u_mem.memory[64] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net449));
 sg13g2_dlygate4sd3_1 hold78 (.A(_0163_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net450));
 sg13g2_dlygate4sd3_1 hold79 (.A(\ppwm_i.u_ppwm.u_mem.memory[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net451));
 sg13g2_dlygate4sd3_1 hold80 (.A(\falu_i.falutop.div_inst.a[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net452));
 sg13g2_dlygate4sd3_1 hold81 (.A(_0340_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net453));
 sg13g2_dlygate4sd3_1 hold82 (.A(\ppwm_i.u_ppwm.u_mem.memory[104] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net454));
 sg13g2_dlygate4sd3_1 hold83 (.A(\ppwm_i.u_ppwm.u_mem.memory[40] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net455));
 sg13g2_dlygate4sd3_1 hold84 (.A(_0140_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net456));
 sg13g2_dlygate4sd3_1 hold85 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net457));
 sg13g2_dlygate4sd3_1 hold86 (.A(_0027_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net458));
 sg13g2_dlygate4sd3_1 hold87 (.A(\falu_i.falutop.i2c_inst.state[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net459));
 sg13g2_dlygate4sd3_1 hold88 (.A(_0220_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net460));
 sg13g2_dlygate4sd3_1 hold89 (.A(\ppwm_i.u_ppwm.u_mem.memory[109] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net461));
 sg13g2_dlygate4sd3_1 hold90 (.A(_0208_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net462));
 sg13g2_dlygate4sd3_1 hold91 (.A(\ppwm_i.u_ppwm.u_mem.memory[70] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net463));
 sg13g2_dlygate4sd3_1 hold92 (.A(_0169_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net464));
 sg13g2_dlygate4sd3_1 hold93 (.A(\falu_i.falutop.div_inst.a[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net465));
 sg13g2_dlygate4sd3_1 hold94 (.A(_0341_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net466));
 sg13g2_dlygate4sd3_1 hold95 (.A(\falu_i.falutop.i2c_inst.op[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net467));
 sg13g2_dlygate4sd3_1 hold96 (.A(_0094_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net468));
 sg13g2_dlygate4sd3_1 hold97 (.A(\ppwm_i.u_ppwm.u_mem.memory[54] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net469));
 sg13g2_dlygate4sd3_1 hold98 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net470));
 sg13g2_dlygate4sd3_1 hold99 (.A(_0028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net471));
 sg13g2_dlygate4sd3_1 hold100 (.A(\ppwm_i.u_ppwm.u_mem.memory[35] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net472));
 sg13g2_dlygate4sd3_1 hold101 (.A(_0135_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net473));
 sg13g2_dlygate4sd3_1 hold102 (.A(\ppwm_i.u_ppwm.u_mem.memory[62] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net474));
 sg13g2_dlygate4sd3_1 hold103 (.A(\falu_i.falutop.div_inst.a[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net475));
 sg13g2_dlygate4sd3_1 hold104 (.A(_0338_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net476));
 sg13g2_dlygate4sd3_1 hold105 (.A(\ppwm_i.u_ppwm.u_mem.memory[22] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net477));
 sg13g2_dlygate4sd3_1 hold106 (.A(_0121_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net478));
 sg13g2_dlygate4sd3_1 hold107 (.A(\falu_i.falutop.div_inst.b1[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net479));
 sg13g2_dlygate4sd3_1 hold108 (.A(_1143_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net480));
 sg13g2_dlygate4sd3_1 hold109 (.A(\ppwm_i.u_ppwm.u_mem.memory[36] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net481));
 sg13g2_dlygate4sd3_1 hold110 (.A(\ppwm_i.u_ppwm.u_mem.memory[72] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net482));
 sg13g2_dlygate4sd3_1 hold111 (.A(\ppwm_i.u_ppwm.u_mem.memory[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net483));
 sg13g2_dlygate4sd3_1 hold112 (.A(_0105_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net484));
 sg13g2_dlygate4sd3_1 hold113 (.A(\falu_i.falutop.div_inst.acc[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net485));
 sg13g2_dlygate4sd3_1 hold114 (.A(_0293_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net486));
 sg13g2_dlygate4sd3_1 hold115 (.A(\falu_i.falutop.div_inst.a[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net487));
 sg13g2_dlygate4sd3_1 hold116 (.A(_0339_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net488));
 sg13g2_dlygate4sd3_1 hold117 (.A(\falu_i.falutop.div_inst.acc[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net489));
 sg13g2_dlygate4sd3_1 hold118 (.A(_0288_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net490));
 sg13g2_dlygate4sd3_1 hold119 (.A(\ppwm_i.u_ppwm.u_mem.memory[63] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net491));
 sg13g2_dlygate4sd3_1 hold120 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net492));
 sg13g2_dlygate4sd3_1 hold121 (.A(_0030_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net493));
 sg13g2_dlygate4sd3_1 hold122 (.A(\falu_i.falutop.div_inst.acc[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net494));
 sg13g2_dlygate4sd3_1 hold123 (.A(_0289_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net495));
 sg13g2_dlygate4sd3_1 hold124 (.A(\ppwm_i.u_ppwm.u_mem.memory[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net496));
 sg13g2_dlygate4sd3_1 hold125 (.A(_0114_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net497));
 sg13g2_dlygate4sd3_1 hold126 (.A(\falu_i.falutop.div_inst.acc[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net498));
 sg13g2_dlygate4sd3_1 hold127 (.A(_0287_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net499));
 sg13g2_dlygate4sd3_1 hold128 (.A(\ppwm_i.u_ppwm.u_mem.memory[101] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net500));
 sg13g2_dlygate4sd3_1 hold129 (.A(_0200_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net501));
 sg13g2_dlygate4sd3_1 hold130 (.A(\ppwm_i.u_ppwm.u_mem.memory[89] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net502));
 sg13g2_dlygate4sd3_1 hold131 (.A(_0189_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net503));
 sg13g2_dlygate4sd3_1 hold132 (.A(\ppwm_i.u_ppwm.u_mem.memory[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net504));
 sg13g2_dlygate4sd3_1 hold133 (.A(_0109_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net505));
 sg13g2_dlygate4sd3_1 hold134 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net506));
 sg13g2_dlygate4sd3_1 hold135 (.A(_0025_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net507));
 sg13g2_dlygate4sd3_1 hold136 (.A(\ppwm_i.u_ppwm.u_mem.memory[26] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net508));
 sg13g2_dlygate4sd3_1 hold137 (.A(_0125_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net509));
 sg13g2_dlygate4sd3_1 hold138 (.A(\ppwm_i.u_ppwm.u_mem.memory[85] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net510));
 sg13g2_dlygate4sd3_1 hold139 (.A(_0185_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net511));
 sg13g2_dlygate4sd3_1 hold140 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net512));
 sg13g2_dlygate4sd3_1 hold141 (.A(_1042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net513));
 sg13g2_dlygate4sd3_1 hold142 (.A(_0218_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net514));
 sg13g2_dlygate4sd3_1 hold143 (.A(\ppwm_i.u_ppwm.u_mem.memory[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net515));
 sg13g2_dlygate4sd3_1 hold144 (.A(\ppwm_i.u_ppwm.u_mem.memory[31] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net516));
 sg13g2_dlygate4sd3_1 hold145 (.A(_0130_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net517));
 sg13g2_dlygate4sd3_1 hold146 (.A(\ppwm_i.u_ppwm.u_mem.memory[87] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net518));
 sg13g2_dlygate4sd3_1 hold147 (.A(_0187_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net519));
 sg13g2_dlygate4sd3_1 hold148 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net520));
 sg13g2_dlygate4sd3_1 hold149 (.A(_0026_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net521));
 sg13g2_dlygate4sd3_1 hold150 (.A(\ppwm_i.u_ppwm.u_mem.memory[65] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net522));
 sg13g2_dlygate4sd3_1 hold151 (.A(\ppwm_i.u_ppwm.u_mem.memory[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net523));
 sg13g2_dlygate4sd3_1 hold152 (.A(_0101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net524));
 sg13g2_dlygate4sd3_1 hold153 (.A(\falu_i.falutop.div_inst.i[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net525));
 sg13g2_dlygate4sd3_1 hold154 (.A(_1139_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net526));
 sg13g2_dlygate4sd3_1 hold155 (.A(_0252_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net527));
 sg13g2_dlygate4sd3_1 hold156 (.A(\ppwm_i.u_ppwm.u_mem.memory[106] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net528));
 sg13g2_dlygate4sd3_1 hold157 (.A(_0205_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net529));
 sg13g2_dlygate4sd3_1 hold158 (.A(\ppwm_i.u_ppwm.u_mem.memory[46] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net530));
 sg13g2_dlygate4sd3_1 hold159 (.A(_0145_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net531));
 sg13g2_dlygate4sd3_1 hold160 (.A(\ppwm_i.u_ppwm.u_mem.memory[96] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net532));
 sg13g2_dlygate4sd3_1 hold161 (.A(_0196_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net533));
 sg13g2_dlygate4sd3_1 hold162 (.A(\ppwm_i.u_ppwm.u_mem.memory[32] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net534));
 sg13g2_dlygate4sd3_1 hold163 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net535));
 sg13g2_dlygate4sd3_1 hold164 (.A(_0033_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net536));
 sg13g2_dlygate4sd3_1 hold165 (.A(\ppwm_i.u_ppwm.u_mem.memory[99] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net537));
 sg13g2_dlygate4sd3_1 hold166 (.A(_0199_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net538));
 sg13g2_dlygate4sd3_1 hold167 (.A(\ppwm_i.u_ppwm.u_mem.memory[102] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net539));
 sg13g2_dlygate4sd3_1 hold168 (.A(\ppwm_i.u_ppwm.u_mem.memory[108] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net540));
 sg13g2_dlygate4sd3_1 hold169 (.A(\ppwm_i.u_ppwm.u_mem.memory[88] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net541));
 sg13g2_dlygate4sd3_1 hold170 (.A(\falu_i.falutop.div_inst.quo[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net542));
 sg13g2_dlygate4sd3_1 hold171 (.A(_0271_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net543));
 sg13g2_dlygate4sd3_1 hold172 (.A(\ppwm_i.u_ppwm.u_mem.memory[86] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net544));
 sg13g2_dlygate4sd3_1 hold173 (.A(\ppwm_i.u_ppwm.u_mem.memory[79] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net545));
 sg13g2_dlygate4sd3_1 hold174 (.A(_0178_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net546));
 sg13g2_dlygate4sd3_1 hold175 (.A(\ppwm_i.u_ppwm.u_mem.memory[33] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net547));
 sg13g2_dlygate4sd3_1 hold176 (.A(_0133_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net548));
 sg13g2_dlygate4sd3_1 hold177 (.A(\falu_i.falutop.div_inst.acc[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net549));
 sg13g2_dlygate4sd3_1 hold178 (.A(_0291_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net550));
 sg13g2_dlygate4sd3_1 hold179 (.A(\ppwm_i.u_ppwm.u_mem.memory[78] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net551));
 sg13g2_dlygate4sd3_1 hold180 (.A(_0177_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net552));
 sg13g2_dlygate4sd3_1 hold181 (.A(\ppwm_i.u_ppwm.global_counter[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net553));
 sg13g2_dlygate4sd3_1 hold182 (.A(_0438_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net554));
 sg13g2_dlygate4sd3_1 hold183 (.A(_0053_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net555));
 sg13g2_dlygate4sd3_1 hold184 (.A(\ppwm_i.u_ppwm.u_mem.memory[95] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net556));
 sg13g2_dlygate4sd3_1 hold185 (.A(\ppwm_i.u_ppwm.u_mem.memory[58] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net557));
 sg13g2_dlygate4sd3_1 hold186 (.A(_0157_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net558));
 sg13g2_dlygate4sd3_1 hold187 (.A(\ppwm_i.u_ppwm.u_mem.memory[110] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net559));
 sg13g2_dlygate4sd3_1 hold188 (.A(\ppwm_i.u_ppwm.u_mem.memory[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net560));
 sg13g2_dlygate4sd3_1 hold189 (.A(_0103_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net561));
 sg13g2_dlygate4sd3_1 hold190 (.A(\ppwm_i.u_ppwm.u_mem.memory[98] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net562));
 sg13g2_dlygate4sd3_1 hold191 (.A(\ppwm_i.u_ppwm.u_mem.memory[77] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net843));
 sg13g2_dlygate4sd3_1 hold192 (.A(\ppwm_i.u_ppwm.u_mem.memory[23] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net844));
 sg13g2_dlygate4sd3_1 hold193 (.A(\ppwm_i.u_ppwm.u_mem.memory[29] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net845));
 sg13g2_dlygate4sd3_1 hold194 (.A(_0129_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net846));
 sg13g2_dlygate4sd3_1 hold195 (.A(\ppwm_i.u_ppwm.u_mem.memory[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net847));
 sg13g2_dlygate4sd3_1 hold196 (.A(\falu_i.falutop.i2c_inst.data_in[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net848));
 sg13g2_dlygate4sd3_1 hold197 (.A(_0228_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net849));
 sg13g2_dlygate4sd3_1 hold198 (.A(\falu_i.falutop.i2c_inst.data_in[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net850));
 sg13g2_dlygate4sd3_1 hold199 (.A(_0234_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net851));
 sg13g2_dlygate4sd3_1 hold200 (.A(\ppwm_i.u_ppwm.u_mem.memory[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net852));
 sg13g2_dlygate4sd3_1 hold201 (.A(_0102_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net853));
 sg13g2_dlygate4sd3_1 hold202 (.A(\ppwm_i.u_ppwm.u_mem.memory[43] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net854));
 sg13g2_dlygate4sd3_1 hold203 (.A(_0142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net855));
 sg13g2_dlygate4sd3_1 hold204 (.A(\falu_i.falutop.div_inst.acc[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net856));
 sg13g2_dlygate4sd3_1 hold205 (.A(_0290_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net857));
 sg13g2_dlygate4sd3_1 hold206 (.A(\falu_i.falutop.i2c_inst.data_in[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net858));
 sg13g2_dlygate4sd3_1 hold207 (.A(_0239_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net859));
 sg13g2_dlygate4sd3_1 hold208 (.A(\ppwm_i.u_ppwm.u_mem.memory[44] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net860));
 sg13g2_dlygate4sd3_1 hold209 (.A(\falu_i.falutop.i2c_inst.data_in[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net861));
 sg13g2_dlygate4sd3_1 hold210 (.A(_0242_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net862));
 sg13g2_dlygate4sd3_1 hold211 (.A(\ppwm_i.u_ppwm.u_pwm.counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net863));
 sg13g2_dlygate4sd3_1 hold212 (.A(_0406_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net864));
 sg13g2_dlygate4sd3_1 hold213 (.A(_0044_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net865));
 sg13g2_dlygate4sd3_1 hold214 (.A(\ppwm_i.u_ppwm.u_mem.memory[59] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net866));
 sg13g2_dlygate4sd3_1 hold215 (.A(\ppwm_i.u_ppwm.u_mem.memory[94] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net867));
 sg13g2_dlygate4sd3_1 hold216 (.A(\ppwm_i.u_ppwm.u_mem.memory[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net868));
 sg13g2_dlygate4sd3_1 hold217 (.A(\falu_i.falutop.i2c_inst.data_in[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net869));
 sg13g2_dlygate4sd3_1 hold218 (.A(_0233_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net870));
 sg13g2_dlygate4sd3_1 hold219 (.A(\falu_i.falutop.i2c_inst.data_in[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net871));
 sg13g2_dlygate4sd3_1 hold220 (.A(_0235_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net872));
 sg13g2_dlygate4sd3_1 hold221 (.A(\falu_i.falutop.i2c_inst.data_in[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net873));
 sg13g2_dlygate4sd3_1 hold222 (.A(_0236_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net874));
 sg13g2_dlygate4sd3_1 hold223 (.A(\ppwm_i.u_ppwm.u_mem.memory[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net875));
 sg13g2_dlygate4sd3_1 hold224 (.A(_0119_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net876));
 sg13g2_dlygate4sd3_1 hold225 (.A(\falu_i.falutop.alu_inst.op[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net877));
 sg13g2_dlygate4sd3_1 hold226 (.A(\ppwm_i.u_ppwm.u_mem.memory[84] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net878));
 sg13g2_dlygate4sd3_1 hold227 (.A(\falu_i.falutop.div_inst.acc[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net879));
 sg13g2_dlygate4sd3_1 hold228 (.A(_1213_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net880));
 sg13g2_dlygate4sd3_1 hold229 (.A(\falu_i.falutop.i2c_inst.data_in[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net881));
 sg13g2_dlygate4sd3_1 hold230 (.A(_0232_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net882));
 sg13g2_dlygate4sd3_1 hold231 (.A(\ppwm_i.u_ppwm.u_mem.programming ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net883));
 sg13g2_dlygate4sd3_1 hold232 (.A(_0907_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net884));
 sg13g2_dlygate4sd3_1 hold233 (.A(\ppwm_i.u_ppwm.u_mem.memory[60] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net885));
 sg13g2_dlygate4sd3_1 hold234 (.A(\ppwm_i.u_ppwm.u_mem.memory[80] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net886));
 sg13g2_dlygate4sd3_1 hold235 (.A(\falu_i.falutop.div_inst.start ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net887));
 sg13g2_dlygate4sd3_1 hold236 (.A(\ppwm_i.u_ppwm.u_mem.memory[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net888));
 sg13g2_dlygate4sd3_1 hold237 (.A(\ppwm_i.u_ppwm.u_mem.memory[67] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net889));
 sg13g2_dlygate4sd3_1 hold238 (.A(_0166_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net890));
 sg13g2_dlygate4sd3_1 hold239 (.A(\falu_i.falutop.div_inst.b[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net891));
 sg13g2_dlygate4sd3_1 hold240 (.A(_0331_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net892));
 sg13g2_dlygate4sd3_1 hold241 (.A(\ppwm_i.u_ppwm.u_mem.memory[45] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net893));
 sg13g2_dlygate4sd3_1 hold242 (.A(\falu_i.falutop.i2c_inst.data_in[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net894));
 sg13g2_dlygate4sd3_1 hold243 (.A(_0241_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net895));
 sg13g2_dlygate4sd3_1 hold244 (.A(\ppwm_i.u_ppwm.u_mem.memory[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net896));
 sg13g2_dlygate4sd3_1 hold245 (.A(\ppwm_i.u_ppwm.u_mem.memory[34] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net897));
 sg13g2_dlygate4sd3_1 hold246 (.A(\ppwm_i.u_ppwm.u_mem.memory[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net898));
 sg13g2_dlygate4sd3_1 hold247 (.A(\falu_i.falutop.i2c_inst.data_in[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net899));
 sg13g2_dlygate4sd3_1 hold248 (.A(_0237_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net900));
 sg13g2_dlygate4sd3_1 hold249 (.A(\falu_i.falutop.i2c_inst.data_in[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net901));
 sg13g2_dlygate4sd3_1 hold250 (.A(_0229_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net902));
 sg13g2_dlygate4sd3_1 hold251 (.A(\ppwm_i.u_ppwm.u_mem.memory[66] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net903));
 sg13g2_dlygate4sd3_1 hold252 (.A(\ppwm_i.u_ppwm.u_mem.memory[68] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net904));
 sg13g2_dlygate4sd3_1 hold253 (.A(\falu_i.falutop.div_inst.val[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net905));
 sg13g2_dlygate4sd3_1 hold254 (.A(\falu_i.falutop.div_inst.a[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net906));
 sg13g2_dlygate4sd3_1 hold255 (.A(_0336_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net907));
 sg13g2_dlygate4sd3_1 hold256 (.A(\falu_i.falutop.i2c_inst.data_in[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net908));
 sg13g2_dlygate4sd3_1 hold257 (.A(_0243_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net909));
 sg13g2_dlygate4sd3_1 hold258 (.A(\falu_i.falutop.div_inst.quo[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net910));
 sg13g2_dlygate4sd3_1 hold259 (.A(_1133_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net911));
 sg13g2_dlygate4sd3_1 hold260 (.A(\falu_i.falutop.i2c_inst.data_in[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net912));
 sg13g2_dlygate4sd3_1 hold261 (.A(_0093_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net913));
 sg13g2_dlygate4sd3_1 hold262 (.A(\ppwm_i.u_ppwm.u_mem.memory[105] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net914));
 sg13g2_dlygate4sd3_1 hold263 (.A(\ppwm_i.u_ppwm.u_mem.memory[52] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net915));
 sg13g2_dlygate4sd3_1 hold264 (.A(_0151_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net916));
 sg13g2_dlygate4sd3_1 hold265 (.A(\falu_i.falutop.div_inst.i[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net917));
 sg13g2_dlygate4sd3_1 hold266 (.A(_1142_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net918));
 sg13g2_dlygate4sd3_1 hold267 (.A(_0253_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net919));
 sg13g2_dlygate4sd3_1 hold268 (.A(\falu_i.falutop.div_inst.b[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net920));
 sg13g2_dlygate4sd3_1 hold269 (.A(_0335_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net921));
 sg13g2_dlygate4sd3_1 hold270 (.A(\ppwm_i.u_ppwm.u_mem.memory[74] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net922));
 sg13g2_dlygate4sd3_1 hold271 (.A(_0173_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net923));
 sg13g2_dlygate4sd3_1 hold272 (.A(\ppwm_i.u_ppwm.u_pwm.cmp_value[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net924));
 sg13g2_dlygate4sd3_1 hold273 (.A(_0032_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net925));
 sg13g2_dlygate4sd3_1 hold274 (.A(\falu_i.falutop.i2c_inst.data_in[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net926));
 sg13g2_dlygate4sd3_1 hold275 (.A(_0240_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net927));
 sg13g2_dlygate4sd3_1 hold276 (.A(\ppwm_i.u_ppwm.u_mem.memory[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net928));
 sg13g2_dlygate4sd3_1 hold277 (.A(_0113_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net929));
 sg13g2_dlygate4sd3_1 hold278 (.A(\ppwm_i.u_ppwm.u_mem.memory[83] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net930));
 sg13g2_dlygate4sd3_1 hold279 (.A(\falu_i.falutop.div_inst.acc[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net931));
 sg13g2_dlygate4sd3_1 hold280 (.A(_0292_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net932));
 sg13g2_dlygate4sd3_1 hold281 (.A(\ppwm_i.u_ppwm.u_mem.memory[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net933));
 sg13g2_dlygate4sd3_1 hold282 (.A(\ppwm_i.u_ppwm.u_mem.data_sync2 ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net934));
 sg13g2_dlygate4sd3_1 hold283 (.A(_1045_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net935));
 sg13g2_dlygate4sd3_1 hold284 (.A(_0219_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net936));
 sg13g2_dlygate4sd3_1 hold285 (.A(\falu_i.falutop.div_inst.val[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net937));
 sg13g2_dlygate4sd3_1 hold286 (.A(\falu_i.falutop.alu_inst.op[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net938));
 sg13g2_dlygate4sd3_1 hold287 (.A(\falu_i.falutop.div_inst.val[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net939));
 sg13g2_dlygate4sd3_1 hold288 (.A(_1147_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net940));
 sg13g2_dlygate4sd3_1 hold289 (.A(_0265_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net941));
 sg13g2_dlygate4sd3_1 hold290 (.A(\ppwm_i.u_ppwm.global_counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net942));
 sg13g2_dlygate4sd3_1 hold291 (.A(_0424_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net943));
 sg13g2_dlygate4sd3_1 hold292 (.A(_0046_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net944));
 sg13g2_dlygate4sd3_1 hold293 (.A(\falu_i.falutop.i2c_inst.data_in[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net945));
 sg13g2_dlygate4sd3_1 hold294 (.A(_0238_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net946));
 sg13g2_dlygate4sd3_1 hold295 (.A(\falu_i.falutop.div_inst.val[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net947));
 sg13g2_dlygate4sd3_1 hold296 (.A(\ppwm_i.u_ppwm.u_mem.memory[81] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net948));
 sg13g2_dlygate4sd3_1 hold297 (.A(\ppwm_i.u_ppwm.u_mem.memory[47] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net949));
 sg13g2_dlygate4sd3_1 hold298 (.A(\ppwm_i.u_ppwm.u_mem.memory[25] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net950));
 sg13g2_dlygate4sd3_1 hold299 (.A(\ppwm_i.u_ppwm.u_mem.memory[111] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net951));
 sg13g2_dlygate4sd3_1 hold300 (.A(\falu_i.falutop.div_inst.a[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net952));
 sg13g2_dlygate4sd3_1 hold301 (.A(_2095_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net953));
 sg13g2_dlygate4sd3_1 hold302 (.A(\ppwm_i.u_ppwm.global_counter[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net954));
 sg13g2_dlygate4sd3_1 hold303 (.A(_0443_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net955));
 sg13g2_dlygate4sd3_1 hold304 (.A(_0056_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net956));
 sg13g2_dlygate4sd3_1 hold305 (.A(\ppwm_i.u_ppwm.u_mem.memory[91] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net957));
 sg13g2_dlygate4sd3_1 hold306 (.A(_0190_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net958));
 sg13g2_dlygate4sd3_1 hold307 (.A(\ppwm_i.u_ppwm.u_mem.memory[28] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net959));
 sg13g2_dlygate4sd3_1 hold308 (.A(_0127_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net960));
 sg13g2_dlygate4sd3_1 hold309 (.A(\ppwm_i.u_ppwm.u_mem.memory[97] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net961));
 sg13g2_dlygate4sd3_1 hold310 (.A(\ppwm_i.u_ppwm.u_mem.memory[69] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net962));
 sg13g2_dlygate4sd3_1 hold311 (.A(\ppwm_i.u_ppwm.u_mem.memory[27] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net963));
 sg13g2_dlygate4sd3_1 hold312 (.A(\falu_i.falutop.alu_inst.op[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net964));
 sg13g2_dlygate4sd3_1 hold313 (.A(\ppwm_i.u_ppwm.u_mem.memory[21] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net965));
 sg13g2_dlygate4sd3_1 hold314 (.A(_0120_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net966));
 sg13g2_dlygate4sd3_1 hold315 (.A(\falu_i.falutop.div_inst.b[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net967));
 sg13g2_dlygate4sd3_1 hold316 (.A(_0332_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net968));
 sg13g2_dlygate4sd3_1 hold317 (.A(\ppwm_i.u_ppwm.u_mem.memory[42] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net969));
 sg13g2_dlygate4sd3_1 hold318 (.A(_0141_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net970));
 sg13g2_dlygate4sd3_1 hold319 (.A(\ppwm_i.u_ppwm.u_mem.data_sync2 ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net971));
 sg13g2_dlygate4sd3_1 hold320 (.A(\falu_i.falutop.i2c_inst.data_in[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net972));
 sg13g2_dlygate4sd3_1 hold321 (.A(_0230_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net973));
 sg13g2_dlygate4sd3_1 hold322 (.A(\ppwm_i.u_ppwm.global_counter[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net974));
 sg13g2_dlygate4sd3_1 hold323 (.A(_0448_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net975));
 sg13g2_dlygate4sd3_1 hold324 (.A(_0059_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net976));
 sg13g2_dlygate4sd3_1 hold325 (.A(\ppwm_i.u_ppwm.u_mem.memory[73] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net977));
 sg13g2_dlygate4sd3_1 hold326 (.A(\falu_i.falutop.div_inst.val[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net978));
 sg13g2_dlygate4sd3_1 hold327 (.A(_0266_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net979));
 sg13g2_dlygate4sd3_1 hold328 (.A(\ppwm_i.u_ppwm.u_ex.state_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net980));
 sg13g2_dlygate4sd3_1 hold329 (.A(_2425_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net981));
 sg13g2_dlygate4sd3_1 hold330 (.A(_0000_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net982));
 sg13g2_dlygate4sd3_1 hold331 (.A(\falu_i.falutop.div_inst.b[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net983));
 sg13g2_dlygate4sd3_1 hold332 (.A(_0334_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net984));
 sg13g2_dlygate4sd3_1 hold333 (.A(\falu_i.falutop.i2c_inst.counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net985));
 sg13g2_dlygate4sd3_1 hold334 (.A(_0349_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net986));
 sg13g2_dlygate4sd3_1 hold335 (.A(_0350_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net987));
 sg13g2_dlygate4sd3_1 hold336 (.A(_0351_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net988));
 sg13g2_dlygate4sd3_1 hold337 (.A(\ppwm_i.u_ppwm.global_counter[17] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net989));
 sg13g2_dlygate4sd3_1 hold338 (.A(_0454_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net990));
 sg13g2_dlygate4sd3_1 hold339 (.A(_0062_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net991));
 sg13g2_dlygate4sd3_1 hold340 (.A(\falu_i.falutop.i2c_inst.data_in[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net992));
 sg13g2_dlygate4sd3_1 hold341 (.A(_0231_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net993));
 sg13g2_dlygate4sd3_1 hold342 (.A(\falu_i.falutop.div_inst.b1[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net994));
 sg13g2_dlygate4sd3_1 hold343 (.A(_1144_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net995));
 sg13g2_dlygate4sd3_1 hold344 (.A(\falu_i.falutop.i2c_inst.sda_o ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net996));
 sg13g2_dlygate4sd3_1 hold345 (.A(_1094_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net997));
 sg13g2_dlygate4sd3_1 hold346 (.A(_0244_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net998));
 sg13g2_dlygate4sd3_1 hold347 (.A(\falu_i.falutop.div_inst.b[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net999));
 sg13g2_dlygate4sd3_1 hold348 (.A(_0333_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1000));
 sg13g2_dlygate4sd3_1 hold349 (.A(\falu_i.falutop.i2c_inst.state[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1001));
 sg13g2_dlygate4sd3_1 hold350 (.A(_2447_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1002));
 sg13g2_dlygate4sd3_1 hold351 (.A(\ppwm_i.u_ppwm.global_counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1003));
 sg13g2_dlygate4sd3_1 hold352 (.A(_0047_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1004));
 sg13g2_dlygate4sd3_1 hold353 (.A(\falu_i.falutop.div_inst.b1[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1005));
 sg13g2_dlygate4sd3_1 hold354 (.A(\falu_i.falutop.i2c_inst.counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1006));
 sg13g2_dlygate4sd3_1 hold355 (.A(_0369_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1007));
 sg13g2_dlygate4sd3_1 hold356 (.A(\ppwm_i.u_ppwm.u_mem.memory[48] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1008));
 sg13g2_dlygate4sd3_1 hold357 (.A(\falu_i.falutop.div_inst.acc[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1009));
 sg13g2_dlygate4sd3_1 hold358 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1010));
 sg13g2_dlygate4sd3_1 hold359 (.A(_1035_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1011));
 sg13g2_dlygate4sd3_1 hold360 (.A(_0216_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1012));
 sg13g2_dlygate4sd3_1 hold361 (.A(\falu_i.falutop.i2c_inst.counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1013));
 sg13g2_dlygate4sd3_1 hold362 (.A(_2437_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1014));
 sg13g2_dlygate4sd3_1 hold363 (.A(\falu_i.falutop.i2c_inst.state[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1015));
 sg13g2_dlygate4sd3_1 hold364 (.A(\falu_i.falutop.i2c_inst.counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1016));
 sg13g2_dlygate4sd3_1 hold365 (.A(_0359_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1017));
 sg13g2_dlygate4sd3_1 hold366 (.A(\falu_i.falutop.i2c_inst.result[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1018));
 sg13g2_dlygate4sd3_1 hold367 (.A(_0307_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1019));
 sg13g2_dlygate4sd3_1 hold368 (.A(\falu_i.falutop.i2c_inst.result[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1020));
 sg13g2_dlygate4sd3_1 hold369 (.A(_0306_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1021));
 sg13g2_dlygate4sd3_1 hold370 (.A(\falu_i.falutop.i2c_inst.result[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1022));
 sg13g2_dlygate4sd3_1 hold371 (.A(_0295_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1023));
 sg13g2_dlygate4sd3_1 hold372 (.A(\ppwm_i.u_ppwm.u_pwm.counter[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1024));
 sg13g2_dlygate4sd3_1 hold373 (.A(_0043_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1025));
 sg13g2_dlygate4sd3_1 hold374 (.A(\falu_i.falutop.i2c_inst.op[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1026));
 sg13g2_dlygate4sd3_1 hold375 (.A(_1137_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1027));
 sg13g2_dlygate4sd3_1 hold376 (.A(\falu_i.falutop.i2c_inst.counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1028));
 sg13g2_dlygate4sd3_1 hold377 (.A(\falu_i.falutop.i2c_inst.result[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1029));
 sg13g2_dlygate4sd3_1 hold378 (.A(_0310_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1030));
 sg13g2_dlygate4sd3_1 hold379 (.A(\ppwm_i.u_ppwm.global_counter[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1031));
 sg13g2_dlygate4sd3_1 hold380 (.A(_0064_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1032));
 sg13g2_dlygate4sd3_1 hold381 (.A(\falu_i.falutop.i2c_inst.result[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1033));
 sg13g2_dlygate4sd3_1 hold382 (.A(_0303_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1034));
 sg13g2_dlygate4sd3_1 hold383 (.A(\falu_i.falutop.i2c_inst.result[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1035));
 sg13g2_dlygate4sd3_1 hold384 (.A(_0308_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1036));
 sg13g2_dlygate4sd3_1 hold385 (.A(\falu_i.falutop.div_inst.val[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1037));
 sg13g2_dlygate4sd3_1 hold386 (.A(_0270_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1038));
 sg13g2_dlygate4sd3_1 hold387 (.A(\ppwm_i.u_ppwm.period_start ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1039));
 sg13g2_dlygate4sd3_1 hold388 (.A(_0002_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1040));
 sg13g2_dlygate4sd3_1 hold389 (.A(\falu_i.falutop.i2c_inst.result[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1041));
 sg13g2_dlygate4sd3_1 hold390 (.A(_0302_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1042));
 sg13g2_dlygate4sd3_1 hold391 (.A(\falu_i.falutop.i2c_inst.counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1043));
 sg13g2_dlygate4sd3_1 hold392 (.A(\falu_i.falutop.i2c_inst.data_in[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1044));
 sg13g2_dlygate4sd3_1 hold393 (.A(\falu_i.falutop.i2c_inst.counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1045));
 sg13g2_dlygate4sd3_1 hold394 (.A(_0343_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1046));
 sg13g2_dlygate4sd3_1 hold395 (.A(\falu_i.falutop.i2c_inst.result[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1047));
 sg13g2_dlygate4sd3_1 hold396 (.A(_0297_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1048));
 sg13g2_dlygate4sd3_1 hold397 (.A(\ppwm_i.u_ppwm.u_pwm.counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1049));
 sg13g2_dlygate4sd3_1 hold398 (.A(_0405_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1050));
 sg13g2_dlygate4sd3_1 hold399 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1051));
 sg13g2_dlygate4sd3_1 hold400 (.A(_1028_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1052));
 sg13g2_dlygate4sd3_1 hold401 (.A(_0214_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1053));
 sg13g2_dlygate4sd3_1 hold402 (.A(\falu_i.falutop.div_inst.b[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1054));
 sg13g2_dlygate4sd3_1 hold403 (.A(_0262_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1055));
 sg13g2_dlygate4sd3_1 hold404 (.A(\falu_i.falutop.div_inst.b1[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1056));
 sg13g2_dlygate4sd3_1 hold405 (.A(\falu_i.falutop.i2c_inst.result[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1057));
 sg13g2_dlygate4sd3_1 hold406 (.A(_0296_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1058));
 sg13g2_dlygate4sd3_1 hold407 (.A(\falu_i.falutop.div_inst.b1[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1059));
 sg13g2_dlygate4sd3_1 hold408 (.A(\ppwm_i.u_ppwm.u_pwm.counter[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1060));
 sg13g2_dlygate4sd3_1 hold409 (.A(_0039_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1061));
 sg13g2_dlygate4sd3_1 hold410 (.A(\falu_i.falutop.i2c_inst.result[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1062));
 sg13g2_dlygate4sd3_1 hold411 (.A(_0305_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1063));
 sg13g2_dlygate4sd3_1 hold412 (.A(\falu_i.falutop.i2c_inst.result[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1064));
 sg13g2_dlygate4sd3_1 hold413 (.A(_0304_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1065));
 sg13g2_dlygate4sd3_1 hold414 (.A(\ppwm_i.u_ppwm.u_pwm.counter[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1066));
 sg13g2_dlygate4sd3_1 hold415 (.A(_0414_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1067));
 sg13g2_dlygate4sd3_1 hold416 (.A(_0040_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1068));
 sg13g2_dlygate4sd3_1 hold417 (.A(\falu_i.falutop.i2c_inst.data_in[19] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1069));
 sg13g2_dlygate4sd3_1 hold418 (.A(\falu_i.falutop.i2c_inst.data_in[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1070));
 sg13g2_dlygate4sd3_1 hold419 (.A(\falu_i.falutop.i2c_inst.result[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1071));
 sg13g2_dlygate4sd3_1 hold420 (.A(_0309_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1072));
 sg13g2_dlygate4sd3_1 hold421 (.A(\falu_i.falutop.data_in[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1073));
 sg13g2_dlygate4sd3_1 hold422 (.A(_2100_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1074));
 sg13g2_dlygate4sd3_1 hold423 (.A(_2101_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1075));
 sg13g2_dlygate4sd3_1 hold424 (.A(\ppwm_i.u_ppwm.global_counter[18] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1076));
 sg13g2_dlygate4sd3_1 hold425 (.A(_0063_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1077));
 sg13g2_dlygate4sd3_1 hold426 (.A(\falu_i.falutop.div_inst.b1[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1078));
 sg13g2_dlygate4sd3_1 hold427 (.A(\falu_i.falutop.div_inst.rem[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1079));
 sg13g2_dlygate4sd3_1 hold428 (.A(_1184_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1080));
 sg13g2_dlygate4sd3_1 hold429 (.A(\falu_i.falutop.div_inst.b[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1081));
 sg13g2_dlygate4sd3_1 hold430 (.A(_0329_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1082));
 sg13g2_dlygate4sd3_1 hold431 (.A(\falu_i.falutop.i2c_inst.result[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1083));
 sg13g2_dlygate4sd3_1 hold432 (.A(\falu_i.falutop.i2c_inst.result[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1084));
 sg13g2_dlygate4sd3_1 hold433 (.A(\falu_i.falutop.div_inst.b1[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1085));
 sg13g2_dlygate4sd3_1 hold434 (.A(\falu_i.falutop.data_in[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1086));
 sg13g2_dlygate4sd3_1 hold435 (.A(_0326_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1087));
 sg13g2_dlygate4sd3_1 hold436 (.A(\falu_i.falutop.i2c_inst.result[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1088));
 sg13g2_dlygate4sd3_1 hold437 (.A(\falu_i.falutop.i2c_inst.result[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1089));
 sg13g2_dlygate4sd3_1 hold438 (.A(\ppwm_i.u_ppwm.u_pwm.counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1090));
 sg13g2_dlygate4sd3_1 hold439 (.A(_0038_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1091));
 sg13g2_dlygate4sd3_1 hold440 (.A(\ppwm_i.u_ppwm.global_counter[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1092));
 sg13g2_dlygate4sd3_1 hold441 (.A(_0437_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1093));
 sg13g2_dlygate4sd3_1 hold442 (.A(\ppwm_i.u_ppwm.u_pwm.counter[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1094));
 sg13g2_dlygate4sd3_1 hold443 (.A(_0042_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1095));
 sg13g2_dlygate4sd3_1 hold444 (.A(\ppwm_i.u_ppwm.global_counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1096));
 sg13g2_dlygate4sd3_1 hold445 (.A(\falu_i.falutop.i2c_inst.counter[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1097));
 sg13g2_dlygate4sd3_1 hold446 (.A(\falu_i.falutop.div_inst.rem[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1098));
 sg13g2_dlygate4sd3_1 hold447 (.A(_0273_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1099));
 sg13g2_dlygate4sd3_1 hold448 (.A(\falu_i.falutop.div_inst.rem[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1100));
 sg13g2_dlygate4sd3_1 hold449 (.A(\falu_i.falutop.data_in[11] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1101));
 sg13g2_dlygate4sd3_1 hold450 (.A(_0324_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1102));
 sg13g2_dlygate4sd3_1 hold451 (.A(\falu_i.falutop.data_in[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1103));
 sg13g2_dlygate4sd3_1 hold452 (.A(_0325_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1104));
 sg13g2_dlygate4sd3_1 hold453 (.A(\falu_i.falutop.data_in[14] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1105));
 sg13g2_dlygate4sd3_1 hold454 (.A(\falu_i.falutop.div_inst.rem[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1106));
 sg13g2_dlygate4sd3_1 hold455 (.A(\ppwm_i.u_ppwm.global_counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1107));
 sg13g2_dlygate4sd3_1 hold456 (.A(_0432_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1108));
 sg13g2_dlygate4sd3_1 hold457 (.A(_0049_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1109));
 sg13g2_dlygate4sd3_1 hold458 (.A(\falu_i.falutop.div_inst.rem[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1110));
 sg13g2_dlygate4sd3_1 hold459 (.A(\ppwm_i.u_ppwm.u_pwm.counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1111));
 sg13g2_dlygate4sd3_1 hold460 (.A(_0401_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1112));
 sg13g2_dlygate4sd3_1 hold461 (.A(_0034_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1113));
 sg13g2_dlygate4sd3_1 hold462 (.A(\falu_i.falutop.data_in[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1114));
 sg13g2_dlygate4sd3_1 hold463 (.A(_0317_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1115));
 sg13g2_dlygate4sd3_1 hold464 (.A(\falu_i.falutop.div_inst.rem[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1116));
 sg13g2_dlygate4sd3_1 hold465 (.A(\ppwm_i.u_ppwm.u_pwm.counter[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1117));
 sg13g2_dlygate4sd3_1 hold466 (.A(_0403_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1118));
 sg13g2_dlygate4sd3_1 hold467 (.A(\falu_i.falutop.div_inst.rem[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1119));
 sg13g2_dlygate4sd3_1 hold468 (.A(\ppwm_i.u_ppwm.global_counter[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1120));
 sg13g2_dlygate4sd3_1 hold469 (.A(_0442_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1121));
 sg13g2_dlygate4sd3_1 hold470 (.A(\falu_i.falutop.data_in[10] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1122));
 sg13g2_dlygate4sd3_1 hold471 (.A(\falu_i.falutop.data_in[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1123));
 sg13g2_dlygate4sd3_1 hold472 (.A(\falu_i.falutop.div_inst.rem[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1124));
 sg13g2_dlygate4sd3_1 hold473 (.A(\ppwm_i.u_ppwm.global_counter[16] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1125));
 sg13g2_dlygate4sd3_1 hold474 (.A(_0453_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1126));
 sg13g2_dlygate4sd3_1 hold475 (.A(\falu_i.falutop.data_in[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1127));
 sg13g2_dlygate4sd3_1 hold476 (.A(_0315_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1128));
 sg13g2_dlygate4sd3_1 hold477 (.A(\ppwm_i.u_ppwm.global_counter[13] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1129));
 sg13g2_dlygate4sd3_1 hold478 (.A(_0447_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1130));
 sg13g2_dlygate4sd3_1 hold479 (.A(\falu_i.falutop.alu_data_in[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1131));
 sg13g2_dlygate4sd3_1 hold480 (.A(\falu_i.falutop.i2c_inst.counter[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1132));
 sg13g2_dlygate4sd3_1 hold481 (.A(\falu_i.falutop.div_inst.val[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1133));
 sg13g2_dlygate4sd3_1 hold482 (.A(\ppwm_i.u_ppwm.global_counter[12] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1134));
 sg13g2_dlygate4sd3_1 hold483 (.A(\falu_i.falutop.data_in[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1135));
 sg13g2_dlygate4sd3_1 hold484 (.A(_0316_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1136));
 sg13g2_dlygate4sd3_1 hold485 (.A(\falu_i.falutop.data_in[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1137));
 sg13g2_dlygate4sd3_1 hold486 (.A(_0320_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1138));
 sg13g2_dlygate4sd3_1 hold487 (.A(\ppwm_i.u_ppwm.global_counter[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1139));
 sg13g2_dlygate4sd3_1 hold488 (.A(_0441_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1140));
 sg13g2_dlygate4sd3_1 hold489 (.A(\falu_i.falutop.data_in[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1141));
 sg13g2_dlygate4sd3_1 hold490 (.A(_0314_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1142));
 sg13g2_dlygate4sd3_1 hold491 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1143));
 sg13g2_dlygate4sd3_1 hold492 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1144));
 sg13g2_dlygate4sd3_1 hold493 (.A(\ppwm_i.u_ppwm.global_counter[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1145));
 sg13g2_dlygate4sd3_1 hold494 (.A(_0434_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1146));
 sg13g2_dlygate4sd3_1 hold495 (.A(_0050_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1147));
 sg13g2_dlygate4sd3_1 hold496 (.A(\falu_i.falutop.data_in[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1148));
 sg13g2_dlygate4sd3_1 hold497 (.A(_0313_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1149));
 sg13g2_dlygate4sd3_1 hold498 (.A(\falu_i.falutop.i2c_inst.counter[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1150));
 sg13g2_dlygate4sd3_1 hold499 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1151));
 sg13g2_dlygate4sd3_1 hold500 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1152));
 sg13g2_dlygate4sd3_1 hold501 (.A(\falu_i.falutop.data_in[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1153));
 sg13g2_dlygate4sd3_1 hold502 (.A(_0318_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1154));
 sg13g2_dlygate4sd3_1 hold503 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1155));
 sg13g2_dlygate4sd3_1 hold504 (.A(_1041_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1156));
 sg13g2_dlygate4sd3_1 hold505 (.A(_0217_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1157));
 sg13g2_dlygate4sd3_1 hold506 (.A(\falu_i.falutop.data_in[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1158));
 sg13g2_dlygate4sd3_1 hold507 (.A(_0321_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1159));
 sg13g2_dlygate4sd3_1 hold508 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1160));
 sg13g2_dlygate4sd3_1 hold509 (.A(_0091_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1161));
 sg13g2_dlygate4sd3_1 hold510 (.A(\ppwm_i.u_ppwm.u_ex.cmp_flag_q ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1162));
 sg13g2_dlygate4sd3_1 hold511 (.A(_0481_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1163));
 sg13g2_dlygate4sd3_1 hold512 (.A(_0066_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1164));
 sg13g2_dlygate4sd3_1 hold513 (.A(\ppwm_i.u_ppwm.pwm_value[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1165));
 sg13g2_dlygate4sd3_1 hold514 (.A(\ppwm_i.u_ppwm.pwm_value[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1166));
 sg13g2_dlygate4sd3_1 hold515 (.A(\ppwm_i.u_ppwm.pwm_value[9] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1167));
 sg13g2_dlygate4sd3_1 hold516 (.A(\ppwm_i.u_ppwm.pc[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1168));
 sg13g2_dlygate4sd3_1 hold517 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1169));
 sg13g2_dlygate4sd3_1 hold518 (.A(_0089_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1170));
 sg13g2_dlygate4sd3_1 hold519 (.A(\ppwm_i.u_ppwm.pwm_value[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1171));
 sg13g2_dlygate4sd3_1 hold520 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1172));
 sg13g2_dlygate4sd3_1 hold521 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[0] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1173));
 sg13g2_dlygate4sd3_1 hold522 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1174));
 sg13g2_dlygate4sd3_1 hold523 (.A(_0087_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1175));
 sg13g2_dlygate4sd3_1 hold524 (.A(\ppwm_i.u_ppwm.pwm_value[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1176));
 sg13g2_dlygate4sd3_1 hold525 (.A(\ppwm_i.u_ppwm.u_pwm.counter[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1177));
 sg13g2_dlygate4sd3_1 hold526 (.A(\falu_i.falutop.data_in[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1178));
 sg13g2_dlygate4sd3_1 hold527 (.A(_0328_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1179));
 sg13g2_dlygate4sd3_1 hold528 (.A(\ppwm_i.u_ppwm.global_counter[15] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1180));
 sg13g2_dlygate4sd3_1 hold529 (.A(\ppwm_i.u_ppwm.pwm_value[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1181));
 sg13g2_dlygate4sd3_1 hold530 (.A(_0076_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1182));
 sg13g2_dlygate4sd3_1 hold531 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[4] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1183));
 sg13g2_dlygate4sd3_1 hold532 (.A(\ppwm_i.u_ppwm.global_counter[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1184));
 sg13g2_dlygate4sd3_1 hold533 (.A(_0436_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1185));
 sg13g2_dlygate4sd3_1 hold534 (.A(\ppwm_i.u_ppwm.u_mem.bit_count[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1186));
 sg13g2_dlygate4sd3_1 hold535 (.A(\ppwm_i.u_ppwm.pwm_value[6] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1187));
 sg13g2_dlygate4sd3_1 hold536 (.A(\ppwm_i.u_ppwm.pwm_value[5] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1188));
 sg13g2_dlygate4sd3_1 hold537 (.A(\ppwm_i.u_ppwm.global_counter[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1189));
 sg13g2_dlygate4sd3_1 hold538 (.A(\ppwm_i.u_ppwm.pwm_value[7] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1190));
 sg13g2_dlygate4sd3_1 hold539 (.A(_0079_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1191));
 sg13g2_dlygate4sd3_1 hold540 (.A(\ppwm_i.u_ppwm.pc[3] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1192));
 sg13g2_dlygate4sd3_1 hold541 (.A(\ppwm_i.u_ppwm.pc[2] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1193));
 sg13g2_dlygate4sd3_1 hold542 (.A(\ppwm_i.u_ppwm.u_ex.reg_value_q[8] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1194));
 sg13g2_dlygate4sd3_1 hold543 (.A(_0090_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1195));
 sg13g2_dlygate4sd3_1 hold544 (.A(\ppwm_i.u_ppwm.pwm_value[1] ),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1196));
 sg13g2_dlygate4sd3_1 hold545 (.A(_0073_),
    .VDD(VPWR),
    .VSS(VGND),
    .X(net1197));
 sg13g2_decap_8 FILLER_0_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_84 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_122 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_168 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_370 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_483 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_539 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_0_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_0_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_0_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_0_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_1_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_1_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_1_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_1_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_86 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_428 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_435 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_550 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_716 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_2_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_2_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_2_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_2_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_585 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_705 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_3_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_733 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_3_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_3_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_3_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_26 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_110 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_137 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_359 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_592 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_4_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_4_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_4_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_4_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_98 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_5_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_5_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_5_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_5_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_19 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_750 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_6_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_6_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_836 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_892 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_899 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_913 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_920 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_6_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_6_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_336 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_567 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_7_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_7_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_7_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_7_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_88 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_515 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_646 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_8_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_8_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_8_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_8_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_522 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_9_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_9_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_9_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_9_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_10 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_50 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_159 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_10_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_10_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_10_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_10_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_322 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_414 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_754 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_11_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_11_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_11_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_11_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_68 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_138 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_280 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_477 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_693 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_759 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_12_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_12_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_12_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_12_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_60 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_139 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_325 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_335 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_355 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_426 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_501 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_736 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_13_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_13_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_13_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_13_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_66 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_167 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_265 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_538 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_641 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_14_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_14_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_14_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_14_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_181 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_220 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_417 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_586 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_674 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_15_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_15_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_15_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_15_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_52 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_56 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_77 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_175 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_263 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_535 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_16_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_16_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_16_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_16_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_314 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_639 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_709 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_719 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_764 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_17_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_834 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_17_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_17_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_17_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_82 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_89 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_374 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_513 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_541 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_548 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_552 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_617 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_18_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_18_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_18_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_18_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_58 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_527 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_773 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_19_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_19_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_19_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_19_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_40 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_42 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_70 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_357 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_382 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_605 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_20_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_20_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_804 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_846 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_20_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_20_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_87 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_160 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_537 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_557 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_21_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_661 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_724 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_726 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_21_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_21_766 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_791 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_805 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_833 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_882 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_21_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_67 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_74 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_97 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_178 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_410 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_571 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_656 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_22_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_22_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_803 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_22_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_22_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_22 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_29 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_36 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_189 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_310 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_312 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_396 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_594 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_601 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_644 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_651 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_23_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_685 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_737 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_744 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_772 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_779 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_807 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_821 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_828 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_849 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_856 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_884 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_891 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_912 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_23_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_23_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_23_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_39 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_46 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_129 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_208 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_219 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_452 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_459 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_528 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_532 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_566 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_24_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_650 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_746 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_760 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_795 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_844 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_24_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_24_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_24_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_48 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_72 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_78 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_150 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_492 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_703 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_728 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_25_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_848 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_855 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_862 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_869 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_876 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_25_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_25_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_25_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_25 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_27 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_51 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_440 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_521 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_26_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_640 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_669 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_681 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_26_842 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_26_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_26_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_80 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_148 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_157 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_207 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_291 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_554 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_570 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_734 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_749 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_27_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_27_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_27_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_889 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_896 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_27_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_28 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_35 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_44 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_83 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_393 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_397 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_563 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_569 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_578 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_606 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_621 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_648 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_730 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_813 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_28_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_28_822 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_28_878 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_903 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_917 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_28_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_194 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_196 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_404 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_468 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_686 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_29_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_29_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_29_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_29_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_16 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_133 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_135 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_163 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_182 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_391 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_451 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_456 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_476 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_534 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_599 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_652 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_662 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_768 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_781 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_30_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_30_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_30_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_30_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_73 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_75 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_180 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_214 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_273 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_318 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_411 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_487 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_591 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_877 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_31_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_31_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_31_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_31_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_53 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_121 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_127 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_162 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_174 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_347 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_425 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_447 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_574 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_630 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_643 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_663 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_670 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_790 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_826 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_854 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_32_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_906 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_32_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_32_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_32_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_32 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_134 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_145 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_152 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_164 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_215 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_224 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_262 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_324 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_341 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_470 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_505 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_507 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_519 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_628 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_642 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_735 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_778 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_798 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_835 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_881 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_33_898 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_33_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_33_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_33_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_8 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_13 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_45 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_57 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_59 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_94 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_228 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_257 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_320 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_500 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_525 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_565 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_608 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_615 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_672 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_694 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_713 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_34_722 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_34_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_34_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_34_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_69 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_115 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_140 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_147 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_149 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_154 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_218 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_226 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_247 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_337 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_344 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_352 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_354 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_395 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_402 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_432 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_514 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_598 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_626 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_738 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_745 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_816 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_35_823 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_910 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_35_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_35_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_35_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_9 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_93 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_107 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_124 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_126 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_239 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_253 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_296 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_303 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_305 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_398 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_409 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_430 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_436 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_443 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_472 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_479 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_484 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_529 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_564 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_579 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_638 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_667 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_680 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_36_700 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_732 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_785 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_843 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_850 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_857 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_36_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_36_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_36_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_61 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_271 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_317 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_330 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_490 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_494 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_556 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_572 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_581 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_633 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_665 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_702 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_758 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_37_771 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_775 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_782 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_831 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_838 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_863 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_870 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_37_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_37_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_37_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_11 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_17 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_24 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_47 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_109 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_116 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_245 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_261 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_268 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_275 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_298 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_331 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_345 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_399 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_419 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_421 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_445 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_512 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_542 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_597 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_612 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_619 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_637 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_654 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_678 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_747 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_752 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_767 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_780 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_789 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_871 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_38_885 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_38_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_38_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_38_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_62 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_91 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_95 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_184 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_191 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_222 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_229 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_284 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_286 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_316 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_323 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_349 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_361 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_363 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_378 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_531 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_549 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_575 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_582 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_636 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_687 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_708 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_712 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_731 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_769 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_840 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_847 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_39_860 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_39_864 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_39_905 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_39_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_37 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_76 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_92 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_99 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_101 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_156 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_166 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_210 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_234 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_241 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_243 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_301 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_315 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_343 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_386 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_416 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_423 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_437 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_454 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_461 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_495 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_499 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_506 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_511 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_518 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_520 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_562 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_593 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_600 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_622 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_629 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_710 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_739 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_756 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_40_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_818 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_825 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_832 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_40_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_40_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_40_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_18 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_20 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_43 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_103 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_114 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_128 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_146 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_153 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_161 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_165 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_201 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_203 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_213 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_233 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_281 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_334 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_353 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_376 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_390 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_408 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_431 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_491 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_498 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_583 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_607 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_614 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_632 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_634 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_649 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_658 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_682 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_689 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_696 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_742 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_757 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_41_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_837 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_41_874 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_927 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_934 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_941 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_948 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_955 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_962 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_969 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_976 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_983 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_990 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_997 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1004 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1011 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_41_1018 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_41_1025 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_85 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_136 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_212 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_216 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_235 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_242 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_249 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_299 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_319 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_342 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_356 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_371 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_384 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_488 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_504 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_524 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_545 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_587 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_664 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_699 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_701 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_720 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_729 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_740 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_751 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_42_761 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_765 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_774 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_786 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_793 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_800 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_810 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_42_820 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_42_853 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_924 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_931 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_938 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_945 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_952 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_959 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_966 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_973 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_980 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_987 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_994 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1001 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1008 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1015 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_42_1022 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_55 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_102 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_117 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_130 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_142 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_176 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_183 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_190 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_192 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_199 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_206 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_236 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_274 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_289 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_302 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_339 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_346 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_350 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_360 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_367 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_380 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_387 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_406 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_438 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_450 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_540 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_547 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_561 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_611 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_624 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_631 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_635 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_647 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_655 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_657 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_762 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_776 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_799 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_806 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_43_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_919 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_926 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_933 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_940 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_947 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_954 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_961 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_968 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_975 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_982 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_989 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_996 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1003 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1010 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_43_1017 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_43_1024 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_43_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_2 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_63 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_65 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_143 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_185 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_187 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_197 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_221 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_225 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_231 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_240 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_260 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_264 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_270 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_272 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_278 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_282 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_306 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_348 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_373 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_375 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_401 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_415 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_422 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_429 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_464 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_471 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_517 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_530 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_536 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_568 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_576 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_603 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_613 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_645 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_671 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_677 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_684 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_691 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_695 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_715 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_717 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_753 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_755 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_44_783 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_44_827 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_44_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_44_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_15 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_30 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_96 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_100 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_105 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_112 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_119 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_132 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_195 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_204 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_238 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_250 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_256 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_267 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_285 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_292 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_294 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_321 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_327 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_377 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_388 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_403 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_442 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_449 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_466 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_473 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_480 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_510 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_523 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_533 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_676 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_787 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_45_797 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_45_867 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_45_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_45_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_4 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_38 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_123 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_171 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_193 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_200 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_217 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_246 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_254 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_313 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_338 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_364 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_366 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_372 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_379 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_385 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_394 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_400 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_407 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_413 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_439 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_446 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_453 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_457 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_486 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_493 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_497 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_544 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_551 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_558 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_573 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_580 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_590 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_595 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_609 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_616 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_623 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_660 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_666 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_673 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_698 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_46_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_46_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_888 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_895 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_902 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_909 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_916 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_923 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_930 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_937 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_944 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_951 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_958 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_965 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_972 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_979 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_986 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_993 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1000 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1007 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1014 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_46_1021 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_46_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_90 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_106 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_113 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_120 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_179 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_186 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_188 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_202 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_209 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_211 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_223 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_232 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_252 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_266 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_328 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_332 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_362 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_381 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_383 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_418 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_433 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_444 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_460 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_467 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_474 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_481 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_508 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_543 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_706 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_743 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_792 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_796 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_802 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_809 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_811 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_817 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_47_829 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_861 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_868 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_875 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_883 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_890 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_897 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_904 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_911 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_918 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_925 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_932 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_939 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_946 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_953 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_960 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_967 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_974 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_981 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_988 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_995 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1002 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1009 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_47_1016 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_47_1023 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_47_1027 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_125 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_155 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_248 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_255 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_259 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_293 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_295 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_300 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_307 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_311 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_369 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_463 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_465 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_526 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_555 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_559 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_620 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_627 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_48_688 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_692 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_707 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_714 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_721 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_723 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_812 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_814 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_851 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_858 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_865 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_872 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_879 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_886 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_893 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_900 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_907 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_914 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_921 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_928 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_935 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_942 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_949 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_956 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_963 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_970 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_977 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_984 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_991 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_998 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1005 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1012 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_48_1019 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_48_1026 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_48_1028 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_0 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_7 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_14 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_21 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_64 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_71 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_79 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_81 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_104 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_111 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_118 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_141 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_151 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_173 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_198 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_205 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_230 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_237 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_244 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_251 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_258 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_269 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_276 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_283 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_290 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_297 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_304 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_309 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_326 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_333 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_340 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_351 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_358 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_365 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_392 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_405 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_412 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_420 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_427 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_434 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_441 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_448 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_455 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_462 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_469 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_475 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_482 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_489 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_496 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_502 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_509 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_516 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_546 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_553 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_560 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_577 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_584 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_588 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_602 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_604 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_618 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_625 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_659 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_668 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_675 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_683 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_690 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_697 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_704 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_711 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_718 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_725 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_727 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_741 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_748 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_763 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_770 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_777 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_784 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_788 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_794 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_801 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_808 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_815 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_819 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_824 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_4 FILLER_49_830 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_839 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_1 FILLER_49_841 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_845 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_852 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_859 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_866 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_873 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_880 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_887 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_894 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_901 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_908 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_915 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_922 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_929 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_936 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_943 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_950 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_957 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_964 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_971 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_978 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_985 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_992 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_999 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1006 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1013 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_decap_8 FILLER_49_1020 (.VDD(VPWR),
    .VSS(VGND));
 sg13g2_fill_2 FILLER_49_1027 (.VDD(VPWR),
    .VSS(VGND));
 assign uio_oe[0] = net8;
 assign uio_oe[1] = net9;
 assign uio_oe[2] = net10;
 assign uio_oe[3] = net11;
 assign uio_oe[4] = net12;
 assign uio_oe[5] = net13;
 assign uio_oe[6] = net14;
 assign uio_oe[7] = net15;
 assign uio_out[0] = net16;
 assign uio_out[1] = net17;
 assign uio_out[2] = net18;
 assign uio_out[3] = net19;
 assign uio_out[4] = net20;
 assign uio_out[5] = net21;
 assign uio_out[6] = net22;
 assign uio_out[7] = net23;
 assign uo_out[1] = net24;
 assign uo_out[2] = net25;
 assign uo_out[3] = net26;
 assign uo_out[5] = net27;
 assign uo_out[6] = net28;
 assign uo_out[7] = net29;
endmodule
