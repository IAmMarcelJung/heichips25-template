* NGSPICE file created from heichips25_tiny_wrapper.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_2 abstract view
.subckt sg13g2_inv_2 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_dlygate4sd3_1 abstract view
.subckt sg13g2_dlygate4sd3_1 A VDD VSS X
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_2 abstract view
.subckt sg13g2_dfrbpq_2 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor2_2 abstract view
.subckt sg13g2_nor2_2 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_2 abstract view
.subckt sg13g2_buf_2 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_2 abstract view
.subckt sg13g2_nand2_2 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_2 abstract view
.subckt sg13g2_nor2b_2 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_and4_1 abstract view
.subckt sg13g2_and4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_inv_4 abstract view
.subckt sg13g2_inv_4 A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_2 abstract view
.subckt sg13g2_nand2b_2 Y B VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_a21o_2 abstract view
.subckt sg13g2_a21o_2 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and3_2 abstract view
.subckt sg13g2_and3_2 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_8 abstract view
.subckt sg13g2_inv_8 Y A VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_2 abstract view
.subckt sg13g2_nor3_2 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

.subckt heichips25_tiny_wrapper VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_39_244 VPWR VGND sg13g2_fill_2
XFILLER_39_222 VPWR VGND sg13g2_decap_8
X_3155_ VGND VPWR net801 _0380_ _0021_ _0381_ sg13g2_a21oi_1
X_3086_ VGND VPWR net800 _2435_ _0003_ _2436_ sg13g2_a21oi_1
XFILLER_36_962 VPWR VGND sg13g2_decap_8
XFILLER_23_601 VPWR VGND sg13g2_fill_2
XFILLER_23_623 VPWR VGND sg13g2_fill_2
XFILLER_23_634 VPWR VGND sg13g2_decap_4
XFILLER_23_667 VPWR VGND sg13g2_fill_1
X_3988_ VGND VPWR net378 _1022_ _0212_ _1023_ sg13g2_a21oi_1
X_2939_ _2293_ net467 VPWR VGND sg13g2_inv_2
X_4609_ _1554_ VPWR _1558_ VGND _1555_ _1556_ sg13g2_o21ai_1
Xhold362 _2437_ VPWR VGND net1014 sg13g2_dlygate4sd3_1
Xhold340 falu_i.falutop.i2c_inst.data_in\[3\] VPWR VGND net992 sg13g2_dlygate4sd3_1
Xhold351 ppwm_i.u_ppwm.global_counter\[2\] VPWR VGND net1003 sg13g2_dlygate4sd3_1
Xhold373 _0043_ VPWR VGND net1025 sg13g2_dlygate4sd3_1
Xhold384 _0308_ VPWR VGND net1036 sg13g2_dlygate4sd3_1
Xhold395 falu_i.falutop.i2c_inst.result\[2\] VPWR VGND net1047 sg13g2_dlygate4sd3_1
Xfanout820 net823 net820 VPWR VGND sg13g2_buf_8
Xfanout842 rst_n net842 VPWR VGND sg13g2_buf_8
Xfanout831 net832 net831 VPWR VGND sg13g2_buf_8
XFILLER_46_748 VPWR VGND sg13g2_fill_1
XFILLER_45_269 VPWR VGND sg13g2_fill_1
XFILLER_27_973 VPWR VGND sg13g2_decap_8
XFILLER_13_100 VPWR VGND sg13g2_fill_2
XFILLER_41_431 VPWR VGND sg13g2_fill_1
XFILLER_41_420 VPWR VGND sg13g2_fill_2
XFILLER_26_85 VPWR VGND sg13g2_fill_2
XFILLER_26_494 VPWR VGND sg13g2_decap_4
XFILLER_42_987 VPWR VGND sg13g2_decap_8
XFILLER_9_126 VPWR VGND sg13g2_decap_8
XFILLER_13_188 VPWR VGND sg13g2_fill_2
XFILLER_10_873 VPWR VGND sg13g2_decap_8
XFILLER_6_899 VPWR VGND sg13g2_decap_8
X_5349__354 VPWR VGND net354 sg13g2_tiehi
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_37_748 VPWR VGND sg13g2_fill_1
XFILLER_36_269 VPWR VGND sg13g2_decap_8
X_4960_ _1903_ net718 _1803_ VPWR VGND sg13g2_nand2_1
XFILLER_18_984 VPWR VGND sg13g2_decap_8
X_3911_ net839 VPWR _0984_ VGND net404 net649 sg13g2_o21ai_1
X_4891_ _1835_ VPWR _1836_ VGND net744 net563 sg13g2_o21ai_1
X_3842_ VGND VPWR _2207_ net641 _0140_ _0949_ sg13g2_a21oi_1
X_5512_ net237 VGND VPWR net543 falu_i.falutop.div_inst.val\[7\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_3773_ net827 VPWR _0915_ VGND net483 net654 sg13g2_o21ai_1
X_5443_ net118 VGND VPWR net393 ppwm_i.u_ppwm.u_mem.memory\[102\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_5374_ net304 VGND VPWR net548 ppwm_i.u_ppwm.u_mem.memory\[33\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_4325_ _1274_ _1276_ _1277_ _1278_ VPWR VGND sg13g2_nor3_1
X_4256_ _1211_ VPWR _0292_ VGND _1098_ _1175_ sg13g2_o21ai_1
X_3207_ _2275_ _0407_ _0411_ _0415_ VPWR VGND sg13g2_nor3_1
X_4187_ _1161_ _1119_ _1120_ VPWR VGND sg13g2_xnor2_1
X_3138_ _2439_ net1007 _0370_ VPWR VGND sg13g2_nor2_1
XFILLER_27_247 VPWR VGND sg13g2_fill_2
XFILLER_24_921 VPWR VGND sg13g2_decap_8
X_3069_ _2422_ _2421_ _2423_ VPWR VGND sg13g2_nor2b_1
XFILLER_24_998 VPWR VGND sg13g2_decap_8
XFILLER_3_803 VPWR VGND sg13g2_decap_4
XFILLER_3_847 VPWR VGND sg13g2_decap_8
XFILLER_2_313 VPWR VGND sg13g2_fill_2
Xhold170 falu_i.falutop.div_inst.quo\[6\] VPWR VGND net542 sg13g2_dlygate4sd3_1
Xhold181 ppwm_i.u_ppwm.global_counter\[8\] VPWR VGND net553 sg13g2_dlygate4sd3_1
Xhold192 ppwm_i.u_ppwm.u_mem.memory\[23\] VPWR VGND net844 sg13g2_dlygate4sd3_1
Xfanout650 net651 net650 VPWR VGND sg13g2_buf_8
Xfanout683 _0386_ net683 VPWR VGND sg13g2_buf_8
Xfanout672 net675 net672 VPWR VGND sg13g2_buf_8
Xfanout661 net663 net661 VPWR VGND sg13g2_buf_8
Xfanout694 net695 net694 VPWR VGND sg13g2_buf_8
XFILLER_18_203 VPWR VGND sg13g2_decap_4
XFILLER_19_737 VPWR VGND sg13g2_decap_8
XFILLER_15_910 VPWR VGND sg13g2_decap_8
XFILLER_42_740 VPWR VGND sg13g2_fill_1
XFILLER_27_792 VPWR VGND sg13g2_fill_2
XFILLER_42_751 VPWR VGND sg13g2_fill_2
XFILLER_15_987 VPWR VGND sg13g2_decap_8
XFILLER_18_1026 VPWR VGND sg13g2_fill_2
XFILLER_41_283 VPWR VGND sg13g2_fill_1
XFILLER_30_979 VPWR VGND sg13g2_decap_8
XFILLER_10_681 VPWR VGND sg13g2_decap_8
XFILLER_6_641 VPWR VGND sg13g2_decap_8
XFILLER_6_696 VPWR VGND sg13g2_fill_1
XFILLER_5_162 VPWR VGND sg13g2_fill_2
X_5090_ _2024_ _2029_ _2030_ VPWR VGND sg13g2_and2_1
X_4110_ falu_i.falutop.div_inst.b1\[5\] falu_i.falutop.div_inst.acc\[5\] _1112_ VPWR
+ VGND sg13g2_nor2b_1
X_5503__269 VPWR VGND net269 sg13g2_tiehi
X_4041_ _1065_ _1059_ _1053_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_556 VPWR VGND sg13g2_fill_2
XFILLER_25_707 VPWR VGND sg13g2_decap_8
X_4943_ VGND VPWR net775 falu_i.falutop.div_inst.rem\[0\] _1887_ falu_i.falutop.div_inst.rem\[1\]
+ sg13g2_a21oi_1
X_4874_ _1819_ _1800_ _1817_ _1818_ VPWR VGND sg13g2_and3_1
XFILLER_21_924 VPWR VGND sg13g2_decap_8
X_3825_ net826 VPWR _0941_ VGND net534 net658 sg13g2_o21ai_1
X_3756_ net807 net375 _0098_ VPWR VGND sg13g2_and2_1
X_3687_ _0840_ _0838_ _0839_ _0849_ VPWR VGND sg13g2_a21o_1
X_5426_ net188 VGND VPWR net511 ppwm_i.u_ppwm.u_mem.memory\[85\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_0_806 VPWR VGND sg13g2_decap_8
X_5357_ net338 VGND VPWR net448 ppwm_i.u_ppwm.u_mem.memory\[16\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_5288_ net121 VGND VPWR net1147 ppwm_i.u_ppwm.global_counter\[5\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
X_4308_ _1259_ _1260_ _1261_ VPWR VGND sg13g2_nor2_2
X_4239_ net542 net605 _1202_ VPWR VGND sg13g2_nor2_1
XFILLER_15_206 VPWR VGND sg13g2_fill_2
XFILLER_28_578 VPWR VGND sg13g2_fill_1
XFILLER_12_902 VPWR VGND sg13g2_decap_8
XFILLER_23_272 VPWR VGND sg13g2_fill_2
XFILLER_24_795 VPWR VGND sg13g2_decap_8
XFILLER_12_979 VPWR VGND sg13g2_decap_8
XFILLER_48_1019 VPWR VGND sg13g2_decap_8
X_5268__160 VPWR VGND net160 sg13g2_tiehi
XFILLER_2_176 VPWR VGND sg13g2_fill_2
XFILLER_19_534 VPWR VGND sg13g2_decap_8
XFILLER_19_556 VPWR VGND sg13g2_decap_4
XFILLER_46_364 VPWR VGND sg13g2_fill_2
XFILLER_34_504 VPWR VGND sg13g2_fill_1
XFILLER_14_283 VPWR VGND sg13g2_decap_4
XFILLER_15_784 VPWR VGND sg13g2_fill_2
XFILLER_30_721 VPWR VGND sg13g2_fill_2
X_3610_ net572 _0774_ _0778_ _0779_ VPWR VGND sg13g2_nor3_1
X_4590_ _1538_ _1537_ _1539_ VPWR VGND sg13g2_xor2_1
X_3541_ _0618_ _0711_ _0712_ _0713_ VPWR VGND sg13g2_nor3_1
XFILLER_7_972 VPWR VGND sg13g2_decap_8
X_3472_ _0646_ VPWR _0647_ VGND _2247_ net596 sg13g2_o21ai_1
X_5211_ VGND VPWR net623 _2124_ _0334_ _2123_ sg13g2_a21oi_1
X_5142_ _2078_ _2079_ _2077_ _2080_ VPWR VGND sg13g2_mux2_1
XFILLER_29_0 VPWR VGND sg13g2_fill_2
X_5073_ _1973_ net773 falu_i.falutop.div_inst.rem\[4\] _2014_ VPWR VGND sg13g2_a21o_1
X_4024_ _1051_ net2 _1050_ VPWR VGND sg13g2_nand2_1
XFILLER_25_559 VPWR VGND sg13g2_fill_2
XFILLER_40_518 VPWR VGND sg13g2_fill_2
XFILLER_12_209 VPWR VGND sg13g2_fill_2
X_4926_ _1851_ _1867_ _1869_ _1870_ VPWR VGND sg13g2_or3_1
X_4857_ _1802_ net752 net727 net768 net712 VPWR VGND sg13g2_a22oi_1
XFILLER_20_264 VPWR VGND sg13g2_fill_1
XFILLER_21_798 VPWR VGND sg13g2_decap_8
X_3808_ VGND VPWR _2218_ net661 _0123_ _0932_ sg13g2_a21oi_1
XFILLER_5_909 VPWR VGND sg13g2_decap_8
X_4788_ _1733_ VPWR _1734_ VGND _1240_ _1314_ sg13g2_o21ai_1
X_3739_ _0887_ _0885_ _0894_ _0896_ VPWR VGND sg13g2_a21o_1
XFILLER_4_419 VPWR VGND sg13g2_decap_8
X_5409_ net234 VGND VPWR _0168_ ppwm_i.u_ppwm.u_mem.memory\[68\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_47_106 VPWR VGND sg13g2_decap_8
X_5380__292 VPWR VGND net292 sg13g2_tiehi
XFILLER_28_386 VPWR VGND sg13g2_decap_8
XFILLER_28_397 VPWR VGND sg13g2_fill_2
XFILLER_43_367 VPWR VGND sg13g2_decap_4
XFILLER_8_703 VPWR VGND sg13g2_fill_1
XFILLER_12_743 VPWR VGND sg13g2_fill_2
XFILLER_4_964 VPWR VGND sg13g2_decap_8
XFILLER_3_496 VPWR VGND sg13g2_fill_1
X_5304__95 VPWR VGND net95 sg13g2_tiehi
XFILLER_19_320 VPWR VGND sg13g2_decap_8
XFILLER_19_342 VPWR VGND sg13g2_decap_4
XFILLER_19_353 VPWR VGND sg13g2_fill_1
XFILLER_34_367 VPWR VGND sg13g2_fill_1
XFILLER_35_879 VPWR VGND sg13g2_decap_8
X_2972_ _2325_ VPWR _2326_ VGND ppwm_i.u_ppwm.u_mem.memory\[36\] _2313_ sg13g2_o21ai_1
X_4711_ _1656_ _1651_ _1658_ VPWR VGND sg13g2_xor2_1
X_4642_ net640 _1589_ _1590_ VPWR VGND sg13g2_nor2_2
X_4573_ _1458_ _1522_ _1523_ VPWR VGND sg13g2_and2_1
X_3524_ _0696_ VPWR _0697_ VGND net584 _0633_ sg13g2_o21ai_1
X_3455_ VPWR _0631_ _0630_ VGND sg13g2_inv_1
X_3386_ ppwm_i.u_ppwm.global_counter\[8\] net782 _0564_ VPWR VGND sg13g2_xor2_1
X_5125_ VGND VPWR _2019_ _2035_ _2064_ _2034_ sg13g2_a21oi_1
X_5056_ _1997_ _1992_ _1995_ VPWR VGND sg13g2_xnor2_1
X_4007_ ppwm_i.u_ppwm.u_mem.bit_count\[4\] ppwm_i.u_ppwm.u_mem.bit_count\[3\] ppwm_i.u_ppwm.u_mem.bit_count\[5\]
+ _1038_ VPWR VGND sg13g2_nand3_1
XFILLER_40_315 VPWR VGND sg13g2_decap_4
X_4909_ _1853_ net727 net751 VPWR VGND sg13g2_nand2_1
X_5289__119 VPWR VGND net119 sg13g2_tiehi
XFILLER_5_717 VPWR VGND sg13g2_fill_2
XFILLER_5_706 VPWR VGND sg13g2_decap_8
XFILLER_1_945 VPWR VGND sg13g2_decap_8
Xhold41 falu_i.falutop.div_inst.b\[1\] VPWR VGND net413 sg13g2_dlygate4sd3_1
Xhold30 ppwm_i.u_ppwm.u_mem.memory\[24\] VPWR VGND net402 sg13g2_dlygate4sd3_1
Xhold52 ppwm_i.u_ppwm.u_mem.memory\[37\] VPWR VGND net424 sg13g2_dlygate4sd3_1
Xhold63 falu_i.falutop.div_inst.quo\[3\] VPWR VGND net435 sg13g2_dlygate4sd3_1
Xhold74 _0206_ VPWR VGND net446 sg13g2_dlygate4sd3_1
Xhold85 ppwm_i.u_ppwm.u_pwm.cmp_value\[3\] VPWR VGND net457 sg13g2_dlygate4sd3_1
XFILLER_17_813 VPWR VGND sg13g2_decap_8
XFILLER_21_1022 VPWR VGND sg13g2_decap_8
Xhold96 _0094_ VPWR VGND net468 sg13g2_dlygate4sd3_1
XFILLER_16_312 VPWR VGND sg13g2_fill_2
XFILLER_43_142 VPWR VGND sg13g2_fill_1
XFILLER_16_378 VPWR VGND sg13g2_fill_2
XFILLER_25_890 VPWR VGND sg13g2_decap_8
XFILLER_31_337 VPWR VGND sg13g2_fill_1
XFILLER_8_522 VPWR VGND sg13g2_decap_8
XFILLER_8_533 VPWR VGND sg13g2_fill_2
XFILLER_8_566 VPWR VGND sg13g2_fill_1
X_3240_ _0435_ net1185 _0051_ VPWR VGND sg13g2_nor2b_1
X_3171_ net810 VPWR _0391_ VGND ppwm_i.u_ppwm.pwm_value\[4\] net683 sg13g2_o21ai_1
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_437 VPWR VGND sg13g2_fill_2
XFILLER_47_481 VPWR VGND sg13g2_decap_8
X_5359__334 VPWR VGND net334 sg13g2_tiehi
XFILLER_23_849 VPWR VGND sg13g2_decap_8
X_2955_ net792 net793 _2309_ VPWR VGND sg13g2_nor2_1
X_2886_ _2240_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] VPWR VGND sg13g2_inv_2
X_4625_ _1074_ VPWR _1574_ VGND _1238_ _1325_ sg13g2_o21ai_1
Xhold511 _0481_ VPWR VGND net1163 sg13g2_dlygate4sd3_1
X_4556_ _1228_ VPWR _1506_ VGND _1230_ _1427_ sg13g2_o21ai_1
Xhold500 ppwm_i.u_ppwm.u_mem.bit_count\[1\] VPWR VGND net1152 sg13g2_dlygate4sd3_1
Xhold533 _0436_ VPWR VGND net1185 sg13g2_dlygate4sd3_1
Xhold522 ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] VPWR VGND net1174 sg13g2_dlygate4sd3_1
Xhold544 ppwm_i.u_ppwm.pwm_value\[1\] VPWR VGND net1196 sg13g2_dlygate4sd3_1
X_3507_ _2272_ net594 _0681_ VPWR VGND sg13g2_nor2_1
X_4487_ VGND VPWR _1291_ _1340_ _1438_ _1337_ sg13g2_a21oi_1
XFILLER_44_1000 VPWR VGND sg13g2_decap_8
X_3438_ VGND VPWR _2255_ _0614_ _0613_ _0611_ sg13g2_a21oi_2
X_3369_ _0546_ VPWR _0547_ VGND _2243_ ppwm_i.u_ppwm.global_counter\[9\] sg13g2_o21ai_1
X_5108_ falu_i.falutop.div_inst.rem\[5\] _2014_ net773 _2048_ VPWR VGND sg13g2_nand3_1
X_5039_ _1788_ _1828_ _1980_ VPWR VGND _1979_ sg13g2_nand3b_1
XFILLER_40_101 VPWR VGND sg13g2_fill_1
XFILLER_14_838 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_4
XFILLER_40_156 VPWR VGND sg13g2_fill_1
XFILLER_31_53 VPWR VGND sg13g2_fill_2
XFILLER_31_75 VPWR VGND sg13g2_fill_1
XFILLER_5_569 VPWR VGND sg13g2_fill_2
Xoutput7 net7 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_45_985 VPWR VGND sg13g2_decap_8
XFILLER_44_473 VPWR VGND sg13g2_fill_1
XFILLER_16_175 VPWR VGND sg13g2_decap_8
XFILLER_31_112 VPWR VGND sg13g2_decap_4
XFILLER_9_853 VPWR VGND sg13g2_decap_8
XFILLER_8_374 VPWR VGND sg13g2_fill_2
X_4410_ VGND VPWR net707 net566 _1362_ _1361_ sg13g2_a21oi_1
X_5390_ net272 VGND VPWR _0149_ ppwm_i.u_ppwm.u_mem.memory\[49\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4341_ _1294_ _2296_ _1292_ VPWR VGND sg13g2_nand2b_1
X_4272_ net760 net730 _1225_ VPWR VGND sg13g2_xor2_1
X_3223_ net942 ppwm_i.u_ppwm.global_counter\[0\] ppwm_i.u_ppwm.period_start _0425_
+ VPWR VGND sg13g2_nand3_1
XFILLER_39_267 VPWR VGND sg13g2_decap_8
XFILLER_11_0 VPWR VGND sg13g2_fill_1
X_3154_ net821 VPWR _0381_ VGND net912 _0380_ sg13g2_o21ai_1
XFILLER_39_278 VPWR VGND sg13g2_fill_1
X_5476__333 VPWR VGND net333 sg13g2_tiehi
X_3085_ net820 VPWR _2436_ VGND net1069 _2435_ sg13g2_o21ai_1
XFILLER_36_941 VPWR VGND sg13g2_decap_8
XFILLER_35_473 VPWR VGND sg13g2_decap_4
X_3987_ net808 VPWR _1023_ VGND net378 net680 sg13g2_o21ai_1
XFILLER_22_178 VPWR VGND sg13g2_fill_2
X_2938_ _2292_ net428 VPWR VGND sg13g2_inv_2
XFILLER_11_1021 VPWR VGND sg13g2_decap_8
X_2869_ VPWR _2223_ net447 VGND sg13g2_inv_1
X_4608_ _1554_ _1555_ _1556_ _1557_ VPWR VGND sg13g2_or3_1
XFILLER_2_528 VPWR VGND sg13g2_decap_4
X_4539_ _1489_ _1429_ _1487_ _1488_ VPWR VGND sg13g2_and3_1
Xhold341 _0231_ VPWR VGND net993 sg13g2_dlygate4sd3_1
Xhold330 _0000_ VPWR VGND net982 sg13g2_dlygate4sd3_1
Xhold352 _0047_ VPWR VGND net1004 sg13g2_dlygate4sd3_1
Xhold385 falu_i.falutop.div_inst.val\[6\] VPWR VGND net1037 sg13g2_dlygate4sd3_1
Xhold396 _0297_ VPWR VGND net1048 sg13g2_dlygate4sd3_1
Xhold363 falu_i.falutop.i2c_inst.state\[0\] VPWR VGND net1015 sg13g2_dlygate4sd3_1
Xhold374 falu_i.falutop.i2c_inst.op\[1\] VPWR VGND net1026 sg13g2_dlygate4sd3_1
Xfanout821 net822 net821 VPWR VGND sg13g2_buf_8
Xfanout832 net833 net832 VPWR VGND sg13g2_buf_2
Xfanout810 net811 net810 VPWR VGND sg13g2_buf_8
XFILLER_19_919 VPWR VGND sg13g2_decap_8
XFILLER_45_204 VPWR VGND sg13g2_fill_2
XFILLER_26_440 VPWR VGND sg13g2_fill_1
XFILLER_27_952 VPWR VGND sg13g2_decap_8
Xclkbuf_3_6__f_clk clknet_0_clk clknet_3_6__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_42_966 VPWR VGND sg13g2_decap_8
XFILLER_13_112 VPWR VGND sg13g2_fill_2
XFILLER_41_498 VPWR VGND sg13g2_decap_4
XFILLER_42_85 VPWR VGND sg13g2_fill_1
XFILLER_10_852 VPWR VGND sg13g2_decap_8
XFILLER_6_878 VPWR VGND sg13g2_decap_8
XFILLER_5_355 VPWR VGND sg13g2_decap_8
XFILLER_3_1008 VPWR VGND sg13g2_decap_8
X_5278__140 VPWR VGND net140 sg13g2_tiehi
XFILLER_18_963 VPWR VGND sg13g2_decap_8
XFILLER_44_270 VPWR VGND sg13g2_fill_2
X_3910_ VGND VPWR _2182_ net678 _0174_ _0983_ sg13g2_a21oi_1
X_4890_ VGND VPWR _2301_ net564 _1835_ _1282_ sg13g2_a21oi_1
XFILLER_17_495 VPWR VGND sg13g2_fill_2
X_3841_ net825 VPWR _0949_ VGND ppwm_i.u_ppwm.u_mem.memory\[41\] net642 sg13g2_o21ai_1
XFILLER_20_605 VPWR VGND sg13g2_decap_8
XFILLER_33_988 VPWR VGND sg13g2_decap_8
XFILLER_32_498 VPWR VGND sg13g2_decap_4
X_3772_ VGND VPWR _2231_ net654 _0105_ _0914_ sg13g2_a21oi_1
X_5511_ net241 VGND VPWR net1038 falu_i.falutop.div_inst.val\[6\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_2
X_5442_ net122 VGND VPWR _0201_ ppwm_i.u_ppwm.u_mem.memory\[101\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_5373_ net306 VGND VPWR _0132_ ppwm_i.u_ppwm.u_mem.memory\[32\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_4324_ _2297_ net747 _1275_ _1277_ VPWR VGND sg13g2_nor3_1
X_4255_ _1211_ net931 net607 VPWR VGND sg13g2_nand2_1
X_3206_ net1066 _0412_ _0414_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1025 VPWR VGND sg13g2_decap_4
X_4186_ VGND VPWR net634 _1159_ _0273_ _1160_ sg13g2_a21oi_1
X_3137_ _0369_ net1006 _0359_ VPWR VGND sg13g2_nand2_2
XFILLER_24_900 VPWR VGND sg13g2_decap_8
X_3068_ _2422_ net419 net821 VPWR VGND sg13g2_nand2_2
XFILLER_11_605 VPWR VGND sg13g2_fill_1
XFILLER_24_977 VPWR VGND sg13g2_decap_8
XFILLER_10_159 VPWR VGND sg13g2_fill_2
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_3_826 VPWR VGND sg13g2_decap_8
Xhold160 ppwm_i.u_ppwm.u_mem.memory\[96\] VPWR VGND net532 sg13g2_dlygate4sd3_1
Xhold171 _0271_ VPWR VGND net543 sg13g2_dlygate4sd3_1
Xhold182 _0438_ VPWR VGND net554 sg13g2_dlygate4sd3_1
Xhold193 ppwm_i.u_ppwm.u_mem.memory\[29\] VPWR VGND net845 sg13g2_dlygate4sd3_1
Xfanout640 _1073_ net640 VPWR VGND sg13g2_buf_8
Xfanout651 net652 net651 VPWR VGND sg13g2_buf_8
Xfanout684 net687 net684 VPWR VGND sg13g2_buf_8
Xfanout673 net675 net673 VPWR VGND sg13g2_buf_8
Xfanout662 net663 net662 VPWR VGND sg13g2_buf_2
Xfanout695 _2311_ net695 VPWR VGND sg13g2_buf_8
XFILLER_42_774 VPWR VGND sg13g2_fill_2
XFILLER_15_966 VPWR VGND sg13g2_decap_8
XFILLER_18_1005 VPWR VGND sg13g2_decap_8
X_5390__272 VPWR VGND net272 sg13g2_tiehi
XFILLER_30_958 VPWR VGND sg13g2_decap_8
XFILLER_10_671 VPWR VGND sg13g2_decap_4
X_5326__49 VPWR VGND net49 sg13g2_tiehi
XFILLER_25_1009 VPWR VGND sg13g2_decap_8
XFILLER_49_351 VPWR VGND sg13g2_decap_8
XFILLER_49_340 VPWR VGND sg13g2_decap_8
X_4040_ VGND VPWR _1059_ _1063_ _0223_ _1064_ sg13g2_a21oi_1
XFILLER_37_502 VPWR VGND sg13g2_fill_2
XFILLER_37_546 VPWR VGND sg13g2_fill_2
XFILLER_18_771 VPWR VGND sg13g2_fill_1
X_4942_ falu_i.falutop.div_inst.rem\[1\] falu_i.falutop.div_inst.rem\[0\] net775 _1886_
+ VPWR VGND sg13g2_nand3_1
XFILLER_21_903 VPWR VGND sg13g2_decap_8
XFILLER_33_763 VPWR VGND sg13g2_fill_1
X_4873_ _1807_ VPWR _1818_ VGND _1814_ _1816_ sg13g2_o21ai_1
XFILLER_33_785 VPWR VGND sg13g2_fill_1
XFILLER_33_796 VPWR VGND sg13g2_fill_2
X_3824_ VGND VPWR _2212_ net657 _0131_ _0940_ sg13g2_a21oi_1
XFILLER_20_479 VPWR VGND sg13g2_decap_8
X_3755_ net807 net374 _0097_ VPWR VGND sg13g2_and2_1
X_3686_ _0848_ _2239_ net600 VPWR VGND sg13g2_xnor2_1
X_5425_ net192 VGND VPWR _0184_ ppwm_i.u_ppwm.u_mem.memory\[84\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_5356_ net340 VGND VPWR _0115_ ppwm_i.u_ppwm.u_mem.memory\[15\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_4307_ _1260_ falu_i.falutop.alu_inst.op\[1\] net877 VPWR VGND sg13g2_nand2_2
X_5287_ net123 VGND VPWR net1109 ppwm_i.u_ppwm.global_counter\[4\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_4238_ VGND VPWR net780 net465 _1201_ _1200_ sg13g2_a21oi_1
XFILLER_28_524 VPWR VGND sg13g2_fill_2
X_4169_ VGND VPWR _2150_ net636 _0267_ _1149_ sg13g2_a21oi_1
XFILLER_24_774 VPWR VGND sg13g2_decap_8
XFILLER_12_958 VPWR VGND sg13g2_decap_8
XFILLER_23_43 VPWR VGND sg13g2_fill_1
XFILLER_7_439 VPWR VGND sg13g2_decap_8
XFILLER_3_667 VPWR VGND sg13g2_decap_8
XFILLER_47_811 VPWR VGND sg13g2_fill_1
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_15_752 VPWR VGND sg13g2_decap_4
XFILLER_31_1024 VPWR VGND sg13g2_decap_4
X_3540_ _0710_ _0709_ _0712_ VPWR VGND sg13g2_nor2b_2
XFILLER_7_951 VPWR VGND sg13g2_decap_8
XFILLER_10_490 VPWR VGND sg13g2_decap_8
X_3471_ _0646_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] net596 VPWR VGND sg13g2_nand2_1
X_5210_ _2124_ falu_i.falutop.data_in\[5\] _2122_ VPWR VGND sg13g2_xnor2_1
X_5247__201 VPWR VGND net201 sg13g2_tiehi
X_5141_ _2078_ VPWR _2079_ VGND _2023_ _2027_ sg13g2_o21ai_1
XFILLER_9_1014 VPWR VGND sg13g2_decap_8
X_5072_ _2010_ _2012_ _1834_ _2013_ VPWR VGND sg13g2_nand3_1
XFILLER_38_811 VPWR VGND sg13g2_fill_2
X_4023_ net1 _1049_ _1050_ VPWR VGND sg13g2_and2_1
X_4925_ VGND VPWR _1865_ _1866_ _1869_ _1852_ sg13g2_a21oi_1
X_4856_ _1801_ net733 net751 VPWR VGND sg13g2_nand2_1
XFILLER_21_755 VPWR VGND sg13g2_fill_1
XFILLER_21_766 VPWR VGND sg13g2_fill_2
X_3807_ net828 VPWR _0932_ VGND ppwm_i.u_ppwm.u_mem.memory\[23\] net661 sg13g2_o21ai_1
X_5369__314 VPWR VGND net314 sg13g2_tiehi
X_5549__259 VPWR VGND net259 sg13g2_tiehi
X_4787_ _1733_ _1240_ _1324_ VPWR VGND sg13g2_nand2_1
XFILLER_20_276 VPWR VGND sg13g2_fill_2
X_3738_ _0887_ _0894_ _0885_ _0895_ VPWR VGND sg13g2_nand3_1
X_3669_ _0824_ _0831_ _0822_ _0833_ VPWR VGND sg13g2_nand3_1
X_5408_ net236 VGND VPWR _0167_ ppwm_i.u_ppwm.u_mem.memory\[67\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
XFILLER_0_604 VPWR VGND sg13g2_decap_8
XFILLER_0_626 VPWR VGND sg13g2_decap_8
X_5339_ net372 VGND VPWR _0098_ ppwm_i.u_ppwm.u_mem.clk_prog_sync3 clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
XFILLER_28_365 VPWR VGND sg13g2_decap_8
XFILLER_43_302 VPWR VGND sg13g2_decap_8
XFILLER_43_346 VPWR VGND sg13g2_decap_4
XFILLER_34_20 VPWR VGND sg13g2_decap_8
X_5491__299 VPWR VGND net299 sg13g2_tiehi
XFILLER_15_1008 VPWR VGND sg13g2_decap_8
XFILLER_4_943 VPWR VGND sg13g2_decap_8
XFILLER_22_508 VPWR VGND sg13g2_fill_1
X_2971_ _2325_ net693 _2205_ net701 _2200_ VPWR VGND sg13g2_a22oi_1
X_4710_ _1657_ _1656_ _1651_ VPWR VGND sg13g2_nand2b_1
XFILLER_15_593 VPWR VGND sg13g2_fill_1
X_4641_ _1259_ _1304_ _1589_ VPWR VGND sg13g2_nor2_1
X_4572_ _1522_ falu_i.falutop.div_inst.val\[2\] _1404_ VPWR VGND sg13g2_nand2_1
X_3523_ _0696_ _0651_ net602 _0631_ net611 VPWR VGND sg13g2_a22oi_1
X_3454_ VGND VPWR _2242_ net598 _0630_ _0629_ sg13g2_a21oi_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_3385_ _2235_ ppwm_i.u_ppwm.global_counter\[9\] _0563_ VPWR VGND sg13g2_nor2_1
X_5124_ _2061_ _2054_ _2063_ VPWR VGND sg13g2_xor2_1
X_5055_ _1992_ _1995_ _1996_ VPWR VGND sg13g2_nor2b_1
X_4006_ VGND VPWR _1034_ net1011 _0216_ _1037_ sg13g2_a21oi_1
XFILLER_26_825 VPWR VGND sg13g2_fill_1
XFILLER_41_806 VPWR VGND sg13g2_fill_2
X_4908_ _1815_ VPWR _1852_ VGND _1807_ _1816_ sg13g2_o21ai_1
X_4839_ net818 VPWR _1785_ VGND net1041 net628 sg13g2_o21ai_1
XFILLER_20_11 VPWR VGND sg13g2_fill_2
XFILLER_1_924 VPWR VGND sg13g2_decap_8
Xhold20 ppwm_i.u_ppwm.u_mem.memory\[103\] VPWR VGND net392 sg13g2_dlygate4sd3_1
Xhold31 _0123_ VPWR VGND net403 sg13g2_dlygate4sd3_1
Xhold53 _0137_ VPWR VGND net425 sg13g2_dlygate4sd3_1
Xhold64 _0282_ VPWR VGND net436 sg13g2_dlygate4sd3_1
Xhold42 _0330_ VPWR VGND net414 sg13g2_dlygate4sd3_1
XFILLER_21_1001 VPWR VGND sg13g2_decap_8
Xhold97 ppwm_i.u_ppwm.u_mem.memory\[54\] VPWR VGND net469 sg13g2_dlygate4sd3_1
Xhold86 _0027_ VPWR VGND net458 sg13g2_dlygate4sd3_1
Xhold75 ppwm_i.u_ppwm.u_mem.memory\[17\] VPWR VGND net447 sg13g2_dlygate4sd3_1
XFILLER_45_30 VPWR VGND sg13g2_fill_2
XFILLER_43_132 VPWR VGND sg13g2_fill_1
XFILLER_17_869 VPWR VGND sg13g2_decap_8
XFILLER_45_96 VPWR VGND sg13g2_decap_4
XFILLER_44_677 VPWR VGND sg13g2_decap_8
XFILLER_43_176 VPWR VGND sg13g2_decap_8
XFILLER_8_545 VPWR VGND sg13g2_fill_2
XFILLER_12_574 VPWR VGND sg13g2_fill_2
XFILLER_4_751 VPWR VGND sg13g2_fill_2
XFILLER_4_784 VPWR VGND sg13g2_decap_8
X_3170_ VGND VPWR _2285_ net683 _0027_ _0390_ sg13g2_a21oi_1
XFILLER_47_460 VPWR VGND sg13g2_fill_2
XFILLER_35_633 VPWR VGND sg13g2_fill_1
XFILLER_23_828 VPWR VGND sg13g2_decap_8
XFILLER_35_677 VPWR VGND sg13g2_fill_2
X_2954_ net788 net700 net786 _2308_ VPWR VGND sg13g2_nand3_1
X_2885_ _2239_ net1183 VPWR VGND sg13g2_inv_2
XFILLER_31_883 VPWR VGND sg13g2_fill_2
X_4624_ _1374_ _1571_ _1572_ _1573_ VPWR VGND sg13g2_nor3_1
Xhold501 falu_i.falutop.data_in\[5\] VPWR VGND net1153 sg13g2_dlygate4sd3_1
X_4555_ _1269_ _1504_ _1505_ VPWR VGND sg13g2_and2_1
Xhold512 _0066_ VPWR VGND net1164 sg13g2_dlygate4sd3_1
Xhold523 _0087_ VPWR VGND net1175 sg13g2_dlygate4sd3_1
Xhold534 ppwm_i.u_ppwm.u_mem.bit_count\[3\] VPWR VGND net1186 sg13g2_dlygate4sd3_1
Xhold545 _0073_ VPWR VGND net1197 sg13g2_dlygate4sd3_1
X_3506_ net586 _0637_ _0680_ VPWR VGND sg13g2_nor2_1
X_4486_ _1434_ _1436_ _1437_ VPWR VGND sg13g2_nor2_1
X_3437_ _0613_ _0612_ net598 VPWR VGND sg13g2_nand2b_1
X_3368_ _0545_ VPWR _0546_ VGND ppwm_i.u_ppwm.pwm_value\[8\] _2267_ sg13g2_o21ai_1
X_5107_ _2014_ net773 falu_i.falutop.div_inst.rem\[5\] _2047_ VPWR VGND sg13g2_a21o_1
XFILLER_46_909 VPWR VGND sg13g2_decap_8
X_3299_ _0480_ VPWR _0481_ VGND _2253_ _0477_ sg13g2_o21ai_1
XFILLER_39_994 VPWR VGND sg13g2_decap_8
X_5038_ _1979_ _1978_ _1879_ VPWR VGND sg13g2_nand2b_1
XFILLER_25_121 VPWR VGND sg13g2_fill_1
XFILLER_41_625 VPWR VGND sg13g2_decap_8
XFILLER_41_614 VPWR VGND sg13g2_decap_8
XFILLER_14_817 VPWR VGND sg13g2_decap_8
XFILLER_41_658 VPWR VGND sg13g2_decap_4
XFILLER_40_113 VPWR VGND sg13g2_fill_2
XFILLER_22_894 VPWR VGND sg13g2_decap_8
XFILLER_5_526 VPWR VGND sg13g2_fill_2
XFILLER_5_548 VPWR VGND sg13g2_decap_4
XFILLER_49_725 VPWR VGND sg13g2_fill_2
XFILLER_0_297 VPWR VGND sg13g2_fill_1
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_29_482 VPWR VGND sg13g2_decap_8
XFILLER_45_964 VPWR VGND sg13g2_decap_8
XFILLER_17_655 VPWR VGND sg13g2_fill_2
XFILLER_17_688 VPWR VGND sg13g2_decap_8
XFILLER_17_699 VPWR VGND sg13g2_fill_1
XFILLER_16_187 VPWR VGND sg13g2_decap_4
XFILLER_31_146 VPWR VGND sg13g2_fill_1
XFILLER_13_894 VPWR VGND sg13g2_decap_8
X_4340_ _2296_ net716 _1293_ VPWR VGND sg13g2_nor2_1
XFILLER_4_592 VPWR VGND sg13g2_fill_1
X_4271_ net732 net757 _1224_ VPWR VGND sg13g2_and2_1
X_3222_ VGND VPWR ppwm_i.u_ppwm.period_start ppwm_i.u_ppwm.global_counter\[0\] _0424_
+ net942 sg13g2_a21oi_1
X_3153_ _2431_ _2446_ _0380_ VPWR VGND sg13g2_nor2_1
X_3084_ _2431_ _2434_ _2435_ VPWR VGND sg13g2_nor2_1
XFILLER_23_603 VPWR VGND sg13g2_fill_1
XFILLER_36_997 VPWR VGND sg13g2_decap_8
XFILLER_23_625 VPWR VGND sg13g2_fill_1
XFILLER_23_658 VPWR VGND sg13g2_decap_8
X_3986_ _1022_ net652 _1021_ VPWR VGND sg13g2_nand2_1
X_5255__185 VPWR VGND net185 sg13g2_tiehi
X_2937_ _2291_ net420 VPWR VGND sg13g2_inv_2
XFILLER_11_1000 VPWR VGND sg13g2_decap_8
X_4607_ _1556_ net756 net741 net762 net737 VPWR VGND sg13g2_a22oi_1
X_2868_ VPWR _2222_ net898 VGND sg13g2_inv_1
X_2799_ VPWR _2153_ net409 VGND sg13g2_inv_1
Xhold320 falu_i.falutop.i2c_inst.data_in\[2\] VPWR VGND net972 sg13g2_dlygate4sd3_1
Xhold342 falu_i.falutop.div_inst.b1\[3\] VPWR VGND net994 sg13g2_dlygate4sd3_1
Xhold353 falu_i.falutop.div_inst.b1\[1\] VPWR VGND net1005 sg13g2_dlygate4sd3_1
X_4538_ _1483_ VPWR _1488_ VGND _1484_ _1486_ sg13g2_o21ai_1
Xhold331 falu_i.falutop.div_inst.b\[5\] VPWR VGND net983 sg13g2_dlygate4sd3_1
Xhold386 _0270_ VPWR VGND net1038 sg13g2_dlygate4sd3_1
X_4469_ _1419_ _1393_ _1420_ VPWR VGND sg13g2_xor2_1
Xhold364 falu_i.falutop.i2c_inst.counter\[4\] VPWR VGND net1016 sg13g2_dlygate4sd3_1
Xfanout800 _2289_ net800 VPWR VGND sg13g2_buf_8
Xhold375 _1137_ VPWR VGND net1027 sg13g2_dlygate4sd3_1
Xfanout822 net823 net822 VPWR VGND sg13g2_buf_8
Xfanout833 net842 net833 VPWR VGND sg13g2_buf_1
Xhold397 ppwm_i.u_ppwm.u_pwm.counter\[2\] VPWR VGND net1049 sg13g2_dlygate4sd3_1
Xfanout811 net814 net811 VPWR VGND sg13g2_buf_8
XFILLER_45_238 VPWR VGND sg13g2_fill_2
XFILLER_27_931 VPWR VGND sg13g2_decap_8
X_5377__298 VPWR VGND net298 sg13g2_tiehi
XFILLER_42_945 VPWR VGND sg13g2_decap_8
XFILLER_41_422 VPWR VGND sg13g2_fill_1
XFILLER_13_102 VPWR VGND sg13g2_fill_1
XFILLER_14_625 VPWR VGND sg13g2_decap_8
XFILLER_41_466 VPWR VGND sg13g2_fill_2
XFILLER_13_146 VPWR VGND sg13g2_decap_4
XFILLER_6_857 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_fill_2
XFILLER_1_551 VPWR VGND sg13g2_fill_2
XFILLER_49_588 VPWR VGND sg13g2_fill_1
XFILLER_49_577 VPWR VGND sg13g2_decap_8
XFILLER_36_205 VPWR VGND sg13g2_decap_4
XFILLER_18_942 VPWR VGND sg13g2_decap_8
XFILLER_44_282 VPWR VGND sg13g2_fill_1
XFILLER_44_260 VPWR VGND sg13g2_decap_4
X_3840_ VGND VPWR _2207_ net653 _0139_ _0948_ sg13g2_a21oi_1
XFILLER_33_967 VPWR VGND sg13g2_decap_8
X_3771_ net824 VPWR _0914_ VGND ppwm_i.u_ppwm.u_mem.memory\[5\] net655 sg13g2_o21ai_1
XFILLER_34_1011 VPWR VGND sg13g2_decap_8
X_5510_ net245 VGND VPWR _0269_ falu_i.falutop.div_inst.val\[5\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_9_695 VPWR VGND sg13g2_decap_8
X_5441_ net126 VGND VPWR net501 ppwm_i.u_ppwm.u_mem.memory\[100\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_2
X_5372_ net308 VGND VPWR _0131_ ppwm_i.u_ppwm.u_mem.memory\[31\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4323_ falu_i.falutop.alu_data_in\[7\] net714 _1276_ VPWR VGND sg13g2_nor2b_1
X_4254_ _1210_ VPWR _0291_ VGND _1098_ _1171_ sg13g2_o21ai_1
XFILLER_41_1004 VPWR VGND sg13g2_decap_8
X_3205_ VGND VPWR _2276_ _0409_ _0039_ _0413_ sg13g2_a21oi_1
X_4185_ net803 VPWR _1160_ VGND net1098 net634 sg13g2_o21ai_1
X_3136_ VGND VPWR net800 _0367_ _0015_ _0368_ sg13g2_a21oi_1
X_3067_ net598 _2420_ _2361_ _2421_ VPWR VGND sg13g2_nand3_1
XFILLER_23_400 VPWR VGND sg13g2_fill_1
XFILLER_24_956 VPWR VGND sg13g2_decap_8
XFILLER_23_488 VPWR VGND sg13g2_decap_8
X_3969_ net841 VPWR _1013_ VGND net454 net673 sg13g2_o21ai_1
Xhold150 ppwm_i.u_ppwm.u_mem.memory\[65\] VPWR VGND net522 sg13g2_dlygate4sd3_1
Xhold161 _0196_ VPWR VGND net533 sg13g2_dlygate4sd3_1
Xhold183 _0053_ VPWR VGND net555 sg13g2_dlygate4sd3_1
Xhold194 _0129_ VPWR VGND net846 sg13g2_dlygate4sd3_1
Xhold172 ppwm_i.u_ppwm.u_mem.memory\[86\] VPWR VGND net544 sg13g2_dlygate4sd3_1
Xfanout630 _1075_ net630 VPWR VGND sg13g2_buf_8
Xfanout641 net642 net641 VPWR VGND sg13g2_buf_8
Xfanout685 net687 net685 VPWR VGND sg13g2_buf_8
Xfanout652 _0908_ net652 VPWR VGND sg13g2_buf_8
Xfanout663 net666 net663 VPWR VGND sg13g2_buf_2
Xfanout674 net675 net674 VPWR VGND sg13g2_buf_2
Xfanout696 net699 net696 VPWR VGND sg13g2_buf_8
XFILLER_46_558 VPWR VGND sg13g2_fill_2
XFILLER_42_720 VPWR VGND sg13g2_decap_8
XFILLER_15_945 VPWR VGND sg13g2_decap_8
XFILLER_27_794 VPWR VGND sg13g2_fill_1
XFILLER_14_455 VPWR VGND sg13g2_fill_2
XFILLER_18_1028 VPWR VGND sg13g2_fill_1
XFILLER_42_786 VPWR VGND sg13g2_decap_8
XFILLER_41_274 VPWR VGND sg13g2_decap_8
XFILLER_30_937 VPWR VGND sg13g2_decap_8
XFILLER_6_687 VPWR VGND sg13g2_fill_1
XFILLER_5_142 VPWR VGND sg13g2_decap_8
XFILLER_45_7 VPWR VGND sg13g2_decap_4
XFILLER_37_558 VPWR VGND sg13g2_fill_1
XFILLER_24_208 VPWR VGND sg13g2_decap_8
X_4941_ _1882_ _1884_ _1834_ _1885_ VPWR VGND sg13g2_nand3_1
XFILLER_24_219 VPWR VGND sg13g2_fill_2
X_4872_ _1807_ _1814_ _1816_ _1817_ VPWR VGND sg13g2_or3_1
X_3823_ net830 VPWR _0940_ VGND net516 net656 sg13g2_o21ai_1
XFILLER_32_274 VPWR VGND sg13g2_decap_8
XFILLER_21_959 VPWR VGND sg13g2_decap_8
XFILLER_20_469 VPWR VGND sg13g2_decap_4
X_3754_ net807 net5 _0096_ VPWR VGND sg13g2_and2_1
X_3685_ _0846_ _0847_ _0085_ VPWR VGND sg13g2_nor2_1
X_5424_ net196 VGND VPWR _0183_ ppwm_i.u_ppwm.u_mem.memory\[83\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
X_5355_ net342 VGND VPWR net497 ppwm_i.u_ppwm.u_mem.memory\[14\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_4306_ _1259_ net772 net771 VPWR VGND sg13g2_nand2_2
X_5286_ net125 VGND VPWR _0048_ ppwm_i.u_ppwm.global_counter\[3\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
X_4237_ net780 _2147_ _1200_ VPWR VGND sg13g2_nor2_1
X_4168_ net818 VPWR _1149_ VGND net947 net636 sg13g2_o21ai_1
X_4099_ VPWR _1102_ _1101_ VGND sg13g2_inv_1
XFILLER_15_208 VPWR VGND sg13g2_fill_1
X_3119_ VGND VPWR net802 _0355_ _0010_ _0356_ sg13g2_a21oi_1
XFILLER_28_569 VPWR VGND sg13g2_decap_8
XFILLER_24_753 VPWR VGND sg13g2_decap_8
XFILLER_11_414 VPWR VGND sg13g2_fill_1
XFILLER_12_937 VPWR VGND sg13g2_decap_8
XFILLER_23_274 VPWR VGND sg13g2_fill_1
XFILLER_23_22 VPWR VGND sg13g2_decap_8
XFILLER_3_646 VPWR VGND sg13g2_fill_2
XFILLER_2_167 VPWR VGND sg13g2_fill_2
XFILLER_2_178 VPWR VGND sg13g2_fill_1
X_5502__271 VPWR VGND net271 sg13g2_tiehi
XFILLER_46_366 VPWR VGND sg13g2_fill_1
XFILLER_15_731 VPWR VGND sg13g2_fill_1
XFILLER_27_591 VPWR VGND sg13g2_decap_8
XFILLER_15_786 VPWR VGND sg13g2_fill_1
XFILLER_14_296 VPWR VGND sg13g2_decap_8
XFILLER_31_1003 VPWR VGND sg13g2_decap_8
XFILLER_7_930 VPWR VGND sg13g2_decap_8
XFILLER_6_495 VPWR VGND sg13g2_decap_8
X_3470_ VPWR VGND _0645_ net799 _0636_ _2251_ _0072_ net573 sg13g2_a221oi_1
XFILLER_43_4 VPWR VGND sg13g2_fill_1
X_5570__64 VPWR VGND net64 sg13g2_tiehi
X_5140_ _2022_ _2021_ _2057_ _2078_ VPWR VGND sg13g2_mux2_1
X_5071_ _2011_ VPWR _2012_ VGND net726 net566 sg13g2_o21ai_1
X_4022_ _2433_ _1048_ _1049_ VPWR VGND sg13g2_nor2_2
X_4924_ _1865_ _1866_ _1852_ _1868_ VPWR VGND sg13g2_nand3_1
X_4855_ _1765_ VPWR _1800_ VGND _1757_ _1766_ sg13g2_o21ai_1
XFILLER_20_211 VPWR VGND sg13g2_fill_2
X_4786_ _1732_ net631 _1731_ VPWR VGND sg13g2_nand2_1
X_3806_ VGND VPWR _2219_ net644 _0122_ _0931_ sg13g2_a21oi_1
X_3737_ _0894_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] net603 VPWR VGND sg13g2_xnor2_1
X_3668_ _0824_ _0822_ _0831_ _0832_ VPWR VGND sg13g2_a21o_1
X_5407_ net238 VGND VPWR net890 ppwm_i.u_ppwm.u_mem.memory\[66\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_3599_ _0768_ _0765_ _0766_ VPWR VGND sg13g2_nand2b_1
X_5338_ net30 VGND VPWR _0097_ ppwm_i.u_ppwm.u_mem.clk_prog_sync2 clknet_leaf_10_clk
+ sg13g2_dfrbpq_1
X_5313__75 VPWR VGND net75 sg13g2_tiehi
X_5269_ net158 VGND VPWR net431 ppwm_i.u_ppwm.u_pwm.cmp_value\[7\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
XFILLER_29_823 VPWR VGND sg13g2_fill_2
XFILLER_34_65 VPWR VGND sg13g2_fill_1
XFILLER_11_244 VPWR VGND sg13g2_fill_2
XFILLER_4_922 VPWR VGND sg13g2_decap_8
XFILLER_4_999 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
X_5463__369 VPWR VGND net369 sg13g2_tiehi
XFILLER_19_300 VPWR VGND sg13g2_decap_4
XFILLER_34_358 VPWR VGND sg13g2_decap_8
X_2970_ net790 VPWR _2324_ VGND ppwm_i.u_ppwm.u_mem.memory\[29\] _2310_ sg13g2_o21ai_1
XFILLER_42_380 VPWR VGND sg13g2_decap_4
X_4640_ _1583_ _1584_ _1588_ _0299_ VPWR VGND sg13g2_nor3_1
X_4571_ net819 VPWR _1521_ VGND net1089 net629 sg13g2_o21ai_1
X_3522_ VPWR _0695_ _0694_ VGND sg13g2_inv_1
XFILLER_6_281 VPWR VGND sg13g2_fill_2
X_3453_ net784 net598 _0629_ VPWR VGND sg13g2_nor2_1
X_3384_ _0562_ _0560_ _0561_ ppwm_i.u_ppwm.global_counter\[7\] _2236_ VPWR VGND sg13g2_a22oi_1
X_5123_ _2054_ _2061_ _2062_ VPWR VGND sg13g2_nor2b_1
X_5405__242 VPWR VGND net242 sg13g2_tiehi
X_5054_ _1995_ _1244_ _1993_ VPWR VGND sg13g2_xnor2_1
X_4005_ _1037_ net807 _1036_ VPWR VGND sg13g2_nand2_1
XFILLER_26_837 VPWR VGND sg13g2_fill_1
XFILLER_38_1009 VPWR VGND sg13g2_decap_8
XFILLER_40_339 VPWR VGND sg13g2_decap_4
X_4907_ _1851_ _1795_ _1850_ VPWR VGND sg13g2_xnor2_1
X_4838_ VPWR VGND net639 _1075_ _1783_ net614 _1784_ _1781_ sg13g2_a221oi_1
XFILLER_14_1020 VPWR VGND sg13g2_decap_8
XFILLER_21_575 VPWR VGND sg13g2_decap_8
X_4769_ _1716_ _1404_ _1646_ VPWR VGND sg13g2_nand2_1
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_fill_1
XFILLER_0_446 VPWR VGND sg13g2_decap_8
XFILLER_49_929 VPWR VGND sg13g2_decap_8
Xhold32 ppwm_i.u_ppwm.u_mem.memory\[76\] VPWR VGND net404 sg13g2_dlygate4sd3_1
XFILLER_0_457 VPWR VGND sg13g2_fill_1
Xhold21 _0202_ VPWR VGND net393 sg13g2_dlygate4sd3_1
Xhold10 _0024_ VPWR VGND net382 sg13g2_dlygate4sd3_1
Xhold43 ppwm_i.u_ppwm.u_mem.memory\[71\] VPWR VGND net415 sg13g2_dlygate4sd3_1
Xhold54 ppwm_i.u_ppwm.u_pwm.cmp_value\[5\] VPWR VGND net426 sg13g2_dlygate4sd3_1
Xhold65 ppwm_i.u_ppwm.u_mem.memory\[61\] VPWR VGND net437 sg13g2_dlygate4sd3_1
Xhold98 ppwm_i.u_ppwm.u_pwm.cmp_value\[4\] VPWR VGND net470 sg13g2_dlygate4sd3_1
Xhold76 _0116_ VPWR VGND net448 sg13g2_dlygate4sd3_1
Xhold87 falu_i.falutop.i2c_inst.state\[1\] VPWR VGND net459 sg13g2_dlygate4sd3_1
XFILLER_16_314 VPWR VGND sg13g2_fill_1
XFILLER_17_848 VPWR VGND sg13g2_decap_8
XFILLER_29_686 VPWR VGND sg13g2_decap_4
XFILLER_44_645 VPWR VGND sg13g2_fill_2
XFILLER_31_306 VPWR VGND sg13g2_fill_1
XFILLER_43_199 VPWR VGND sg13g2_decap_8
XFILLER_40_851 VPWR VGND sg13g2_decap_8
XFILLER_8_502 VPWR VGND sg13g2_decap_4
XFILLER_40_895 VPWR VGND sg13g2_fill_2
X_5387__278 VPWR VGND net278 sg13g2_tiehi
XFILLER_4_741 VPWR VGND sg13g2_fill_1
XFILLER_3_240 VPWR VGND sg13g2_decap_8
XFILLER_6_1018 VPWR VGND sg13g2_decap_8
XFILLER_48_984 VPWR VGND sg13g2_decap_8
XFILLER_22_306 VPWR VGND sg13g2_fill_2
XFILLER_23_807 VPWR VGND sg13g2_decap_8
XFILLER_37_1020 VPWR VGND sg13g2_decap_8
X_2953_ _2307_ net791 net793 VPWR VGND sg13g2_nand2_1
XFILLER_16_881 VPWR VGND sg13g2_decap_8
X_2884_ _2238_ net1174 VPWR VGND sg13g2_inv_2
XFILLER_31_895 VPWR VGND sg13g2_decap_4
X_4623_ _1570_ _1239_ _1572_ VPWR VGND sg13g2_nor2b_1
X_5288__121 VPWR VGND net121 sg13g2_tiehi
Xhold502 _0318_ VPWR VGND net1154 sg13g2_dlygate4sd3_1
X_4554_ _1264_ _1268_ _1225_ _1504_ VPWR VGND sg13g2_nand3_1
Xhold524 ppwm_i.u_ppwm.pwm_value\[8\] VPWR VGND net1176 sg13g2_dlygate4sd3_1
Xhold535 ppwm_i.u_ppwm.pwm_value\[6\] VPWR VGND net1187 sg13g2_dlygate4sd3_1
Xhold513 ppwm_i.u_ppwm.pwm_value\[0\] VPWR VGND net1165 sg13g2_dlygate4sd3_1
X_3505_ VPWR VGND _0622_ _0675_ _0678_ _0627_ _0679_ net571 sg13g2_a221oi_1
X_4485_ _1436_ net615 _1435_ VPWR VGND sg13g2_nand2_1
X_3436_ _2345_ _2360_ _0612_ VPWR VGND sg13g2_nor2_1
X_3367_ _0544_ VPWR _0545_ VGND _0533_ _0543_ sg13g2_o21ai_1
X_5106_ _2043_ _2045_ _1834_ _2046_ VPWR VGND sg13g2_nand3_1
X_3298_ VGND VPWR _2253_ net793 _0480_ _0479_ sg13g2_a21oi_1
XFILLER_39_973 VPWR VGND sg13g2_decap_8
X_5037_ _1920_ _1964_ _1978_ VPWR VGND sg13g2_nor2_1
XFILLER_22_873 VPWR VGND sg13g2_decap_8
XFILLER_1_700 VPWR VGND sg13g2_fill_1
XFILLER_1_744 VPWR VGND sg13g2_decap_8
XFILLER_49_704 VPWR VGND sg13g2_decap_8
XFILLER_49_748 VPWR VGND sg13g2_fill_2
XFILLER_36_409 VPWR VGND sg13g2_fill_2
XFILLER_29_461 VPWR VGND sg13g2_decap_8
XFILLER_45_943 VPWR VGND sg13g2_decap_8
XFILLER_44_464 VPWR VGND sg13g2_decap_8
X_5534__112 VPWR VGND net112 sg13g2_tiehi
XFILLER_32_637 VPWR VGND sg13g2_fill_1
XFILLER_9_811 VPWR VGND sg13g2_fill_2
XFILLER_13_873 VPWR VGND sg13g2_decap_8
XFILLER_9_888 VPWR VGND sg13g2_decap_8
XFILLER_8_376 VPWR VGND sg13g2_fill_1
XFILLER_28_1008 VPWR VGND sg13g2_decap_8
X_4270_ VPWR _1223_ _1222_ VGND sg13g2_inv_1
X_3221_ net795 _0423_ _0045_ VPWR VGND sg13g2_nor2_1
X_3152_ VGND VPWR net800 _0378_ _0020_ _0379_ sg13g2_a21oi_1
X_3083_ _2434_ _2432_ _2433_ VPWR VGND sg13g2_nand2_2
XFILLER_36_976 VPWR VGND sg13g2_decap_8
XFILLER_22_147 VPWR VGND sg13g2_decap_8
X_3985_ _1021_ net934 _0906_ VPWR VGND sg13g2_nand2_2
X_2936_ VPWR _2290_ net485 VGND sg13g2_inv_1
X_2867_ VPWR _2221_ net875 VGND sg13g2_inv_1
XFILLER_30_180 VPWR VGND sg13g2_fill_2
X_4606_ net741 net737 net762 net756 _1555_ VPWR VGND sg13g2_and4_1
Xhold310 ppwm_i.u_ppwm.u_mem.memory\[69\] VPWR VGND net962 sg13g2_dlygate4sd3_1
X_2798_ VPWR _2152_ net910 VGND sg13g2_inv_1
Xhold343 _1144_ VPWR VGND net995 sg13g2_dlygate4sd3_1
X_4537_ _1483_ _1484_ _1486_ _1487_ VPWR VGND sg13g2_or3_1
Xhold332 _0334_ VPWR VGND net984 sg13g2_dlygate4sd3_1
Xhold321 _0230_ VPWR VGND net973 sg13g2_dlygate4sd3_1
X_4468_ _1418_ _1417_ _1419_ VPWR VGND sg13g2_xor2_1
Xhold376 falu_i.falutop.i2c_inst.counter\[1\] VPWR VGND net1028 sg13g2_dlygate4sd3_1
Xhold365 _0359_ VPWR VGND net1017 sg13g2_dlygate4sd3_1
Xhold354 falu_i.falutop.i2c_inst.counter\[2\] VPWR VGND net1006 sg13g2_dlygate4sd3_1
Xhold387 ppwm_i.u_ppwm.period_start VPWR VGND net1039 sg13g2_dlygate4sd3_1
Xfanout834 net835 net834 VPWR VGND sg13g2_buf_8
X_3419_ VPWR VGND _2246_ _0596_ ppwm_i.u_ppwm.global_counter\[16\] _2245_ _0597_ ppwm_i.u_ppwm.global_counter\[17\]
+ sg13g2_a221oi_1
Xhold398 _0405_ VPWR VGND net1050 sg13g2_dlygate4sd3_1
Xfanout801 _2289_ net801 VPWR VGND sg13g2_buf_1
Xfanout823 rst_n net823 VPWR VGND sg13g2_buf_8
Xfanout812 net814 net812 VPWR VGND sg13g2_buf_8
X_4399_ VGND VPWR _1229_ _1252_ _1351_ _1251_ sg13g2_a21oi_1
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_26_44 VPWR VGND sg13g2_decap_8
XFILLER_27_987 VPWR VGND sg13g2_decap_8
XFILLER_42_924 VPWR VGND sg13g2_decap_8
XFILLER_41_412 VPWR VGND sg13g2_fill_2
XFILLER_41_401 VPWR VGND sg13g2_fill_1
XFILLER_14_659 VPWR VGND sg13g2_decap_8
XFILLER_6_803 VPWR VGND sg13g2_decap_8
XFILLER_6_836 VPWR VGND sg13g2_decap_8
XFILLER_6_814 VPWR VGND sg13g2_fill_1
XFILLER_10_887 VPWR VGND sg13g2_decap_8
X_5564__116 VPWR VGND net116 sg13g2_tiehi
XFILLER_18_921 VPWR VGND sg13g2_decap_8
XFILLER_36_239 VPWR VGND sg13g2_decap_4
XFILLER_44_250 VPWR VGND sg13g2_fill_1
XFILLER_44_272 VPWR VGND sg13g2_fill_1
XFILLER_18_998 VPWR VGND sg13g2_decap_8
XFILLER_33_946 VPWR VGND sg13g2_decap_8
XFILLER_32_445 VPWR VGND sg13g2_fill_2
X_3770_ VGND VPWR _2232_ net641 _0104_ _0913_ sg13g2_a21oi_1
XFILLER_41_990 VPWR VGND sg13g2_decap_8
X_5440_ net130 VGND VPWR net538 ppwm_i.u_ppwm.u_mem.memory\[99\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_5371_ net310 VGND VPWR net517 ppwm_i.u_ppwm.u_mem.memory\[30\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_4322_ net714 net705 _1275_ VPWR VGND sg13g2_nor2_1
X_4253_ _1210_ net549 net607 VPWR VGND sg13g2_nand2_1
X_3204_ net809 VPWR _0413_ VGND _0407_ _0411_ sg13g2_o21ai_1
X_4184_ _1158_ VPWR _1159_ VGND net498 net568 sg13g2_o21ai_1
X_3135_ net816 VPWR _0368_ VGND net858 _0367_ sg13g2_o21ai_1
X_3066_ net585 net608 _2420_ VPWR VGND sg13g2_nor2_1
XFILLER_24_935 VPWR VGND sg13g2_decap_8
XFILLER_23_434 VPWR VGND sg13g2_fill_1
XFILLER_11_629 VPWR VGND sg13g2_decap_8
X_3968_ VGND VPWR _2162_ net648 _0203_ _1012_ sg13g2_a21oi_1
X_2919_ _2273_ net1024 VPWR VGND sg13g2_inv_2
X_3899_ net839 VPWR _0978_ VGND ppwm_i.u_ppwm.u_mem.memory\[69\] net676 sg13g2_o21ai_1
XFILLER_12_68 VPWR VGND sg13g2_fill_1
X_5569_ net72 VGND VPWR net1179 falu_i.falutop.alu_data_in\[15\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
Xhold162 ppwm_i.u_ppwm.u_mem.memory\[32\] VPWR VGND net534 sg13g2_dlygate4sd3_1
Xhold140 ppwm_i.u_ppwm.u_mem.bit_count\[6\] VPWR VGND net512 sg13g2_dlygate4sd3_1
Xhold151 ppwm_i.u_ppwm.u_mem.memory\[1\] VPWR VGND net523 sg13g2_dlygate4sd3_1
Xhold173 ppwm_i.u_ppwm.u_mem.memory\[79\] VPWR VGND net545 sg13g2_dlygate4sd3_1
Xhold184 ppwm_i.u_ppwm.u_mem.memory\[95\] VPWR VGND net556 sg13g2_dlygate4sd3_1
Xhold195 ppwm_i.u_ppwm.u_mem.memory\[5\] VPWR VGND net847 sg13g2_dlygate4sd3_1
Xfanout642 net645 net642 VPWR VGND sg13g2_buf_8
Xfanout631 _1306_ net631 VPWR VGND sg13g2_buf_8
Xfanout620 net621 net620 VPWR VGND sg13g2_buf_1
Xfanout664 net665 net664 VPWR VGND sg13g2_buf_8
Xfanout675 net679 net675 VPWR VGND sg13g2_buf_8
Xfanout653 net655 net653 VPWR VGND sg13g2_buf_8
Xfanout686 net687 net686 VPWR VGND sg13g2_buf_2
Xfanout697 net698 net697 VPWR VGND sg13g2_buf_8
XFILLER_27_762 VPWR VGND sg13g2_decap_4
XFILLER_15_924 VPWR VGND sg13g2_decap_8
XFILLER_42_765 VPWR VGND sg13g2_fill_1
XFILLER_41_242 VPWR VGND sg13g2_decap_8
XFILLER_41_231 VPWR VGND sg13g2_fill_2
X_5531__137 VPWR VGND net137 sg13g2_tiehi
XFILLER_2_883 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_4
X_5577__307 VPWR VGND net307 sg13g2_tiehi
XFILLER_18_762 VPWR VGND sg13g2_decap_8
X_4940_ _1883_ VPWR _1884_ VGND net740 net564 sg13g2_o21ai_1
XFILLER_18_795 VPWR VGND sg13g2_decap_8
X_4871_ VGND VPWR _1812_ _1813_ _1816_ _1808_ sg13g2_a21oi_1
X_3822_ VGND VPWR _2213_ net664 _0130_ _0939_ sg13g2_a21oi_1
XFILLER_20_415 VPWR VGND sg13g2_fill_1
XFILLER_21_938 VPWR VGND sg13g2_decap_8
XFILLER_33_798 VPWR VGND sg13g2_fill_1
X_3753_ VGND VPWR _2292_ net686 _0095_ _0905_ sg13g2_a21oi_1
X_5573__40 VPWR VGND net40 sg13g2_tiehi
X_3684_ net822 VPWR _0847_ VGND net1151 _0813_ sg13g2_o21ai_1
X_5423_ net200 VGND VPWR _0182_ ppwm_i.u_ppwm.u_mem.memory\[82\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_5354_ net344 VGND VPWR net929 ppwm_i.u_ppwm.u_mem.memory\[13\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_5325__51 VPWR VGND net51 sg13g2_tiehi
X_4305_ VGND VPWR _1258_ _1256_ _1218_ sg13g2_or2_1
X_5285_ net127 VGND VPWR net1004 ppwm_i.u_ppwm.global_counter\[2\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_4236_ VGND VPWR net606 _1198_ _0284_ _1199_ sg13g2_a21oi_1
X_4167_ VGND VPWR _2151_ net637 _0266_ _1148_ sg13g2_a21oi_1
X_3118_ net804 VPWR _0356_ VGND net850 _0355_ sg13g2_o21ai_1
X_4098_ _1101_ _1099_ _1100_ VPWR VGND sg13g2_nand2_2
XFILLER_28_559 VPWR VGND sg13g2_decap_4
X_3049_ VPWR VGND _2402_ net787 _2401_ _2398_ _2403_ _2400_ sg13g2_a221oi_1
XFILLER_24_732 VPWR VGND sg13g2_decap_8
X_5415__222 VPWR VGND net222 sg13g2_tiehi
XFILLER_12_916 VPWR VGND sg13g2_decap_8
XFILLER_8_909 VPWR VGND sg13g2_decap_8
XFILLER_11_459 VPWR VGND sg13g2_fill_2
XFILLER_20_993 VPWR VGND sg13g2_decap_8
XFILLER_3_603 VPWR VGND sg13g2_fill_1
XFILLER_3_4 VPWR VGND sg13g2_decap_8
X_5422__204 VPWR VGND net204 sg13g2_tiehi
XFILLER_47_802 VPWR VGND sg13g2_decap_8
X_5576__351 VPWR VGND net351 sg13g2_tiehi
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_27_570 VPWR VGND sg13g2_decap_8
XFILLER_34_518 VPWR VGND sg13g2_fill_2
XFILLER_34_529 VPWR VGND sg13g2_fill_1
XFILLER_9_14 VPWR VGND sg13g2_decap_8
XFILLER_9_58 VPWR VGND sg13g2_fill_1
XFILLER_30_768 VPWR VGND sg13g2_fill_1
XFILLER_11_993 VPWR VGND sg13g2_decap_8
XFILLER_7_986 VPWR VGND sg13g2_decap_8
XFILLER_6_452 VPWR VGND sg13g2_decap_8
XFILLER_6_474 VPWR VGND sg13g2_fill_1
X_5070_ VGND VPWR _2303_ net566 _2011_ _1282_ sg13g2_a21oi_1
X_4021_ falu_i.falutop.i2c_inst.state\[0\] net459 _1048_ VPWR VGND sg13g2_nor2b_2
XFILLER_37_334 VPWR VGND sg13g2_fill_2
X_5397__258 VPWR VGND net258 sg13g2_tiehi
X_4923_ _1867_ _1852_ _1865_ _1866_ VPWR VGND sg13g2_and3_1
XFILLER_33_551 VPWR VGND sg13g2_fill_2
X_4854_ _1799_ _1791_ _1797_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_223 VPWR VGND sg13g2_fill_2
XFILLER_21_724 VPWR VGND sg13g2_fill_2
X_4785_ VGND VPWR net632 net565 _1731_ _1730_ sg13g2_a21oi_1
X_3805_ net828 VPWR _0931_ VGND net844 net644 sg13g2_o21ai_1
X_3736_ _0892_ _0893_ _0090_ VPWR VGND sg13g2_nor2_1
XFILLER_20_278 VPWR VGND sg13g2_fill_1
X_3667_ VPWR _0831_ _0830_ VGND sg13g2_inv_1
X_5406_ net240 VGND VPWR _0165_ ppwm_i.u_ppwm.u_mem.memory\[65\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_3598_ _0767_ _0766_ _0765_ VPWR VGND sg13g2_nand2b_1
X_5337_ net31 VGND VPWR _0096_ ppwm_i.u_ppwm.u_mem.clk_prog_sync1 clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_5268_ net160 VGND VPWR net493 ppwm_i.u_ppwm.u_pwm.cmp_value\[6\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_4219_ net399 net606 _1187_ VPWR VGND sg13g2_nor2_1
X_5298__101 VPWR VGND net101 sg13g2_tiehi
X_5199_ VGND VPWR net624 _2115_ _0331_ _2113_ sg13g2_a21oi_1
XFILLER_28_323 VPWR VGND sg13g2_decap_8
XFILLER_44_827 VPWR VGND sg13g2_fill_2
XFILLER_43_326 VPWR VGND sg13g2_decap_8
XFILLER_18_89 VPWR VGND sg13g2_fill_2
XFILLER_12_702 VPWR VGND sg13g2_fill_2
XFILLER_12_713 VPWR VGND sg13g2_decap_8
XFILLER_24_562 VPWR VGND sg13g2_decap_4
XFILLER_8_717 VPWR VGND sg13g2_decap_4
XFILLER_4_901 VPWR VGND sg13g2_decap_8
X_5537__84 VPWR VGND net84 sg13g2_tiehi
XFILLER_4_978 VPWR VGND sg13g2_decap_8
XFILLER_38_109 VPWR VGND sg13g2_decap_8
XFILLER_35_816 VPWR VGND sg13g2_decap_8
XFILLER_46_186 VPWR VGND sg13g2_decap_8
XFILLER_34_326 VPWR VGND sg13g2_decap_8
XFILLER_15_540 VPWR VGND sg13g2_fill_2
XFILLER_15_551 VPWR VGND sg13g2_fill_1
X_4570_ VPWR VGND net616 _1519_ _1461_ _1261_ _1520_ _1410_ sg13g2_a221oi_1
X_3521_ _0694_ net602 net612 VPWR VGND sg13g2_nand2_2
X_3452_ net602 _0621_ _0628_ VPWR VGND sg13g2_nor2_1
X_3383_ _0561_ _2269_ ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] _2268_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\]
+ VPWR VGND sg13g2_a22oi_1
X_5122_ _2060_ _2055_ _2061_ VPWR VGND sg13g2_xor2_1
XFILLER_27_0 VPWR VGND sg13g2_decap_4
X_5053_ net724 net705 _1244_ _1994_ VPWR VGND sg13g2_nor3_1
XFILLER_38_654 VPWR VGND sg13g2_decap_4
X_4004_ ppwm_i.u_ppwm.u_mem.bit_count\[3\] _1030_ net1010 _1036_ VPWR VGND sg13g2_nand3_1
X_5449__91 VPWR VGND net91 sg13g2_tiehi
XFILLER_1_92 VPWR VGND sg13g2_decap_8
XFILLER_26_816 VPWR VGND sg13g2_decap_8
X_4906_ _1850_ _1844_ _1848_ VPWR VGND sg13g2_xnor2_1
X_4837_ _1783_ falu_i.falutop.div_inst.val\[7\] _1782_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_598 VPWR VGND sg13g2_fill_1
X_4768_ _1714_ VPWR _1715_ VGND _1663_ _1664_ sg13g2_o21ai_1
X_3719_ _0876_ _0877_ net575 _0878_ VPWR VGND sg13g2_nand3_1
X_4699_ VGND VPWR net937 _1644_ _1647_ _1074_ sg13g2_a21oi_1
XFILLER_49_908 VPWR VGND sg13g2_decap_8
XFILLER_0_425 VPWR VGND sg13g2_decap_8
XFILLER_1_959 VPWR VGND sg13g2_decap_8
X_5265__166 VPWR VGND net166 sg13g2_tiehi
Xhold11 ppwm_i.u_ppwm.u_mem.memory\[75\] VPWR VGND net383 sg13g2_dlygate4sd3_1
XFILLER_0_469 VPWR VGND sg13g2_decap_8
Xhold22 ppwm_i.u_ppwm.u_mem.memory\[56\] VPWR VGND net394 sg13g2_dlygate4sd3_1
Xhold44 _0170_ VPWR VGND net416 sg13g2_dlygate4sd3_1
Xhold55 _0029_ VPWR VGND net427 sg13g2_dlygate4sd3_1
Xhold33 falu_i.falutop.div_inst.quo\[4\] VPWR VGND net405 sg13g2_dlygate4sd3_1
Xhold66 _0160_ VPWR VGND net438 sg13g2_dlygate4sd3_1
Xhold77 ppwm_i.u_ppwm.u_mem.memory\[64\] VPWR VGND net449 sg13g2_dlygate4sd3_1
Xhold99 _0028_ VPWR VGND net471 sg13g2_dlygate4sd3_1
Xhold88 _0220_ VPWR VGND net460 sg13g2_dlygate4sd3_1
XFILLER_44_613 VPWR VGND sg13g2_fill_1
XFILLER_17_827 VPWR VGND sg13g2_decap_8
XFILLER_43_123 VPWR VGND sg13g2_decap_8
XFILLER_12_521 VPWR VGND sg13g2_fill_2
XFILLER_31_318 VPWR VGND sg13g2_fill_2
XFILLER_12_543 VPWR VGND sg13g2_decap_4
XFILLER_24_392 VPWR VGND sg13g2_fill_1
XFILLER_3_296 VPWR VGND sg13g2_decap_8
XFILLER_0_981 VPWR VGND sg13g2_decap_8
XFILLER_48_963 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_fill_1
XFILLER_19_153 VPWR VGND sg13g2_decap_8
XFILLER_16_860 VPWR VGND sg13g2_decap_8
X_5461__42 VPWR VGND net42 sg13g2_tiehi
X_2952_ net791 net793 _2306_ VPWR VGND sg13g2_and2_1
XFILLER_31_830 VPWR VGND sg13g2_fill_2
X_2883_ _2237_ net1172 VPWR VGND sg13g2_inv_2
XFILLER_31_885 VPWR VGND sg13g2_fill_1
X_4622_ _1224_ _1239_ _1507_ _1571_ VPWR VGND sg13g2_nor3_1
X_4553_ _1502_ _1501_ _1499_ _1503_ VPWR VGND sg13g2_a21o_1
Xhold525 ppwm_i.u_ppwm.u_pwm.counter\[7\] VPWR VGND net1177 sg13g2_dlygate4sd3_1
X_3504_ _0647_ _0677_ net610 _0678_ VPWR VGND sg13g2_mux2_1
Xhold536 ppwm_i.u_ppwm.pwm_value\[5\] VPWR VGND net1188 sg13g2_dlygate4sd3_1
X_4484_ _1379_ VPWR _1435_ VGND _1431_ _1433_ sg13g2_o21ai_1
Xhold503 ppwm_i.u_ppwm.u_mem.bit_count\[5\] VPWR VGND net1155 sg13g2_dlygate4sd3_1
Xhold514 ppwm_i.u_ppwm.pwm_value\[3\] VPWR VGND net1166 sg13g2_dlygate4sd3_1
X_3435_ net579 VPWR _0611_ VGND _0609_ net589 sg13g2_o21ai_1
X_3366_ _0544_ _2268_ ppwm_i.u_ppwm.pwm_value\[7\] _2267_ ppwm_i.u_ppwm.pwm_value\[8\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_44_1014 VPWR VGND sg13g2_decap_8
X_3297_ VGND VPWR _0479_ _0478_ _2329_ sg13g2_or2_1
X_5105_ _2044_ VPWR _2045_ VGND net722 net564 sg13g2_o21ai_1
XFILLER_39_952 VPWR VGND sg13g2_decap_8
X_5036_ VGND VPWR _1972_ _1976_ _0306_ _1977_ sg13g2_a21oi_1
XFILLER_26_602 VPWR VGND sg13g2_decap_8
XFILLER_41_649 VPWR VGND sg13g2_fill_1
XFILLER_22_852 VPWR VGND sg13g2_decap_8
XFILLER_5_528 VPWR VGND sg13g2_fill_1
XFILLER_5_506 VPWR VGND sg13g2_fill_2
XFILLER_0_211 VPWR VGND sg13g2_decap_8
XFILLER_49_727 VPWR VGND sg13g2_fill_1
XFILLER_48_259 VPWR VGND sg13g2_fill_1
XFILLER_48_248 VPWR VGND sg13g2_decap_8
XFILLER_45_922 VPWR VGND sg13g2_decap_8
XFILLER_17_613 VPWR VGND sg13g2_fill_2
XFILLER_17_635 VPWR VGND sg13g2_decap_4
XFILLER_45_999 VPWR VGND sg13g2_decap_8
XFILLER_17_657 VPWR VGND sg13g2_fill_1
XFILLER_13_852 VPWR VGND sg13g2_decap_8
XFILLER_9_867 VPWR VGND sg13g2_decap_8
X_3220_ _0423_ net1039 net1096 VPWR VGND sg13g2_xnor2_1
X_3151_ net820 VPWR _0379_ VGND net1070 _0378_ sg13g2_o21ai_1
X_3082_ net1001 falu_i.falutop.i2c_inst.state\[0\] _2433_ VPWR VGND sg13g2_nor2b_2
XFILLER_35_432 VPWR VGND sg13g2_decap_8
XFILLER_36_955 VPWR VGND sg13g2_decap_8
XFILLER_35_443 VPWR VGND sg13g2_fill_2
X_5552__235 VPWR VGND net235 sg13g2_tiehi
XFILLER_23_616 VPWR VGND sg13g2_decap_8
X_3984_ VGND VPWR _2156_ net646 _0211_ _1020_ sg13g2_a21oi_1
X_2935_ _2289_ net3 VPWR VGND sg13g2_inv_2
X_2866_ VPWR _2220_ net965 VGND sg13g2_inv_1
X_4605_ _1554_ net732 net767 VPWR VGND sg13g2_nand2_1
Xhold300 falu_i.falutop.div_inst.a\[7\] VPWR VGND net952 sg13g2_dlygate4sd3_1
X_2797_ VPWR _2151_ net399 VGND sg13g2_inv_1
Xhold311 ppwm_i.u_ppwm.u_mem.memory\[27\] VPWR VGND net963 sg13g2_dlygate4sd3_1
Xhold322 ppwm_i.u_ppwm.global_counter\[14\] VPWR VGND net974 sg13g2_dlygate4sd3_1
X_4536_ _1486_ net756 net745 net762 net741 VPWR VGND sg13g2_a22oi_1
Xhold333 falu_i.falutop.i2c_inst.counter\[3\] VPWR VGND net985 sg13g2_dlygate4sd3_1
Xhold344 falu_i.falutop.i2c_inst.sda_o VPWR VGND net996 sg13g2_dlygate4sd3_1
Xhold377 falu_i.falutop.i2c_inst.result\[15\] VPWR VGND net1029 sg13g2_dlygate4sd3_1
X_4467_ _1418_ net740 net721 VPWR VGND sg13g2_nand2_1
Xhold366 falu_i.falutop.i2c_inst.result\[12\] VPWR VGND net1018 sg13g2_dlygate4sd3_1
Xhold355 _0369_ VPWR VGND net1007 sg13g2_dlygate4sd3_1
X_3418_ VPWR VGND ppwm_i.u_ppwm.pwm_value\[5\] _0595_ _2262_ ppwm_i.u_ppwm.pwm_value\[6\]
+ _0596_ _2261_ sg13g2_a221oi_1
Xfanout813 net814 net813 VPWR VGND sg13g2_buf_1
X_4398_ _1249_ VPWR _1350_ VGND net632 _1247_ sg13g2_o21ai_1
Xfanout802 _2289_ net802 VPWR VGND sg13g2_buf_8
Xhold399 ppwm_i.u_ppwm.u_mem.bit_count\[2\] VPWR VGND net1051 sg13g2_dlygate4sd3_1
Xfanout824 net832 net824 VPWR VGND sg13g2_buf_8
Xhold388 _0002_ VPWR VGND net1040 sg13g2_dlygate4sd3_1
X_3349_ VPWR VGND _2237_ _0526_ ppwm_i.u_ppwm.pwm_value\[6\] _2236_ _0527_ ppwm_i.u_ppwm.pwm_value\[7\]
+ sg13g2_a221oi_1
Xfanout835 net842 net835 VPWR VGND sg13g2_buf_8
X_5019_ _1960_ _1934_ _1961_ VPWR VGND sg13g2_nor2b_1
XFILLER_27_966 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_decap_8
XFILLER_10_866 VPWR VGND sg13g2_decap_8
XFILLER_49_502 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_decap_8
XFILLER_18_900 VPWR VGND sg13g2_decap_8
XFILLER_29_281 VPWR VGND sg13g2_fill_2
XFILLER_44_240 VPWR VGND sg13g2_fill_2
XFILLER_18_977 VPWR VGND sg13g2_decap_8
X_5370_ net312 VGND VPWR net846 ppwm_i.u_ppwm.u_mem.memory\[29\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_5582__239 VPWR VGND net239 sg13g2_tiehi
XFILLER_5_881 VPWR VGND sg13g2_decap_8
X_4321_ _1274_ net632 _1247_ _1273_ VPWR VGND sg13g2_and3_1
X_4252_ _1209_ VPWR _0290_ VGND _1098_ _1167_ sg13g2_o21ai_1
X_3203_ _0407_ _0411_ _0412_ VPWR VGND sg13g2_nor2_1
X_4183_ _1158_ net568 _1157_ VPWR VGND sg13g2_nand2_1
X_3134_ _2434_ _0360_ _0367_ VPWR VGND sg13g2_nor2_1
XFILLER_27_207 VPWR VGND sg13g2_fill_2
X_3065_ net608 _2419_ VPWR VGND sg13g2_inv_4
XFILLER_35_240 VPWR VGND sg13g2_decap_8
XFILLER_24_914 VPWR VGND sg13g2_decap_8
XFILLER_36_785 VPWR VGND sg13g2_fill_2
X_3967_ net838 VPWR _1012_ VGND net454 net648 sg13g2_o21ai_1
X_2918_ _2272_ net1003 VPWR VGND sg13g2_inv_2
X_3898_ VGND VPWR _2187_ net649 _0168_ _0977_ sg13g2_a21oi_1
XFILLER_12_25 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_30_clk clknet_3_7__leaf_clk clknet_leaf_30_clk VPWR VGND sg13g2_buf_8
X_2849_ VPWR _2203_ net530 VGND sg13g2_inv_1
X_5568_ net80 VGND VPWR _0327_ falu_i.falutop.alu_data_in\[14\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
X_4519_ _1467_ net721 _1468_ _1469_ VPWR VGND sg13g2_a21o_1
Xhold141 _1042_ VPWR VGND net513 sg13g2_dlygate4sd3_1
Xhold130 ppwm_i.u_ppwm.u_mem.memory\[89\] VPWR VGND net502 sg13g2_dlygate4sd3_1
Xhold152 _0101_ VPWR VGND net524 sg13g2_dlygate4sd3_1
Xhold174 _0178_ VPWR VGND net546 sg13g2_dlygate4sd3_1
Xhold163 ppwm_i.u_ppwm.u_pwm.cmp_value\[9\] VPWR VGND net535 sg13g2_dlygate4sd3_1
Xhold185 ppwm_i.u_ppwm.u_mem.memory\[58\] VPWR VGND net557 sg13g2_dlygate4sd3_1
X_5499_ net277 VGND VPWR _0258_ falu_i.falutop.div_inst.b1\[3\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
Xfanout610 _2389_ net610 VPWR VGND sg13g2_buf_8
X_5524__178 VPWR VGND net178 sg13g2_tiehi
Xfanout632 _1242_ net632 VPWR VGND sg13g2_buf_8
Xfanout621 _1136_ net621 VPWR VGND sg13g2_buf_8
Xhold196 falu_i.falutop.i2c_inst.data_in\[0\] VPWR VGND net848 sg13g2_dlygate4sd3_1
Xfanout676 net678 net676 VPWR VGND sg13g2_buf_8
Xfanout665 net666 net665 VPWR VGND sg13g2_buf_8
Xfanout643 net645 net643 VPWR VGND sg13g2_buf_8
Xfanout654 net655 net654 VPWR VGND sg13g2_buf_1
Xfanout698 net699 net698 VPWR VGND sg13g2_buf_8
Xfanout687 _0902_ net687 VPWR VGND sg13g2_buf_8
XFILLER_39_590 VPWR VGND sg13g2_decap_4
XFILLER_18_218 VPWR VGND sg13g2_decap_4
XFILLER_18_229 VPWR VGND sg13g2_fill_1
XFILLER_15_903 VPWR VGND sg13g2_decap_8
XFILLER_27_785 VPWR VGND sg13g2_fill_2
XFILLER_18_1019 VPWR VGND sg13g2_decap_8
XFILLER_14_457 VPWR VGND sg13g2_fill_1
XFILLER_6_612 VPWR VGND sg13g2_fill_2
XFILLER_6_601 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_21_clk clknet_3_6__leaf_clk clknet_leaf_21_clk VPWR VGND sg13g2_buf_8
XFILLER_6_634 VPWR VGND sg13g2_decap_8
X_5466__357 VPWR VGND net357 sg13g2_tiehi
XFILLER_2_862 VPWR VGND sg13g2_decap_8
XFILLER_49_365 VPWR VGND sg13g2_fill_2
X_5473__339 VPWR VGND net339 sg13g2_tiehi
XFILLER_33_722 VPWR VGND sg13g2_decap_4
X_4870_ _1812_ _1813_ _1808_ _1815_ VPWR VGND sg13g2_nand3_1
X_3821_ net830 VPWR _0939_ VGND ppwm_i.u_ppwm.u_mem.memory\[30\] net664 sg13g2_o21ai_1
XFILLER_21_917 VPWR VGND sg13g2_decap_8
XFILLER_20_427 VPWR VGND sg13g2_decap_4
X_3752_ falu_i.falutop.i2c_inst.data_in\[19\] net686 _0905_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_12_clk clknet_3_2__leaf_clk clknet_leaf_12_clk VPWR VGND sg13g2_buf_8
X_3683_ VGND VPWR net575 _0842_ _0846_ _0845_ sg13g2_a21oi_1
X_5422_ net204 VGND VPWR net418 ppwm_i.u_ppwm.u_mem.memory\[81\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_5353_ net346 VGND VPWR _0112_ ppwm_i.u_ppwm.u_mem.memory\[12\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_4304_ _1257_ _1218_ _1256_ VPWR VGND sg13g2_nand2_1
X_5284_ net129 VGND VPWR net944 ppwm_i.u_ppwm.global_counter\[1\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_4235_ net432 net605 _1199_ VPWR VGND sg13g2_nor2_1
X_4166_ net817 VPWR _1148_ VGND net978 net637 sg13g2_o21ai_1
X_3117_ _0344_ net987 _0355_ VPWR VGND sg13g2_nor2_1
X_4097_ net413 net1081 net967 net891 _1100_ VPWR VGND sg13g2_nor4_1
XFILLER_24_711 VPWR VGND sg13g2_decap_8
X_3048_ VPWR VGND _2228_ net790 net689 _2233_ _2402_ net696 sg13g2_a221oi_1
XFILLER_36_593 VPWR VGND sg13g2_fill_1
XFILLER_24_788 VPWR VGND sg13g2_decap_8
X_4999_ _1941_ _1936_ _1940_ VPWR VGND sg13g2_nand2_1
XFILLER_20_972 VPWR VGND sg13g2_decap_8
XFILLER_2_125 VPWR VGND sg13g2_fill_1
XFILLER_48_21 VPWR VGND sg13g2_fill_1
XFILLER_24_1012 VPWR VGND sg13g2_decap_8
XFILLER_46_313 VPWR VGND sg13g2_fill_2
XFILLER_19_527 VPWR VGND sg13g2_decap_8
XFILLER_19_549 VPWR VGND sg13g2_decap_8
XFILLER_46_379 VPWR VGND sg13g2_fill_1
X_5275__146 VPWR VGND net146 sg13g2_tiehi
XFILLER_14_265 VPWR VGND sg13g2_decap_8
XFILLER_15_777 VPWR VGND sg13g2_decap_8
XFILLER_30_714 VPWR VGND sg13g2_decap_8
XFILLER_14_276 VPWR VGND sg13g2_decap_8
XFILLER_11_972 VPWR VGND sg13g2_decap_8
XFILLER_7_965 VPWR VGND sg13g2_decap_8
XFILLER_9_1028 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk clknet_leaf_1_clk VPWR VGND sg13g2_buf_8
X_4020_ net459 _1047_ _0220_ VPWR VGND sg13g2_nor2_1
XFILLER_49_173 VPWR VGND sg13g2_decap_8
XFILLER_49_151 VPWR VGND sg13g2_decap_4
XFILLER_37_346 VPWR VGND sg13g2_fill_1
X_4922_ _1856_ VPWR _1866_ VGND _1862_ _1864_ sg13g2_o21ai_1
X_4853_ _1791_ _1797_ _1798_ VPWR VGND sg13g2_nor2_1
X_4784_ net632 _1667_ _1729_ _1730_ VPWR VGND sg13g2_nor3_1
X_3804_ VGND VPWR _2219_ net661 _0121_ _0930_ sg13g2_a21oi_1
X_3735_ net822 VPWR _0893_ VGND net783 _0813_ sg13g2_o21ai_1
X_5405_ net242 VGND VPWR _0164_ ppwm_i.u_ppwm.u_mem.memory\[64\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_3666_ _0830_ _2241_ net602 VPWR VGND sg13g2_xnor2_1
X_3597_ VGND VPWR net1187 net601 _0766_ _0750_ sg13g2_a21oi_1
XFILLER_47_1023 VPWR VGND sg13g2_decap_4
XFILLER_0_618 VPWR VGND sg13g2_fill_2
X_5336_ net32 VGND VPWR net429 falu_i.falutop.i2c_inst.op\[3\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_5267_ net162 VGND VPWR net427 ppwm_i.u_ppwm.u_pwm.cmp_value\[5\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_4218_ VGND VPWR net779 falu_i.falutop.div_inst.a\[0\] _1186_ _1185_ sg13g2_a21oi_1
XFILLER_18_24 VPWR VGND sg13g2_fill_2
X_5198_ _2114_ falu_i.falutop.data_in\[2\] _2115_ VPWR VGND sg13g2_xor2_1
XFILLER_28_302 VPWR VGND sg13g2_fill_1
X_4149_ VGND VPWR _2153_ _1140_ _0254_ net778 sg13g2_a21oi_1
XFILLER_44_817 VPWR VGND sg13g2_fill_1
XFILLER_28_379 VPWR VGND sg13g2_decap_8
XFILLER_34_45 VPWR VGND sg13g2_fill_2
XFILLER_11_246 VPWR VGND sg13g2_fill_1
Xclkload0 clknet_3_3__leaf_clk clkload0/X VPWR VGND sg13g2_buf_8
XFILLER_4_957 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_decap_4
XFILLER_19_313 VPWR VGND sg13g2_decap_8
XFILLER_19_346 VPWR VGND sg13g2_fill_1
XFILLER_34_316 VPWR VGND sg13g2_decap_4
XFILLER_34_338 VPWR VGND sg13g2_fill_2
XFILLER_42_371 VPWR VGND sg13g2_fill_2
XFILLER_30_588 VPWR VGND sg13g2_fill_2
XFILLER_30_599 VPWR VGND sg13g2_decap_4
XFILLER_11_791 VPWR VGND sg13g2_decap_4
X_3520_ _0692_ VPWR _0693_ VGND _0688_ _0691_ sg13g2_o21ai_1
XFILLER_7_762 VPWR VGND sg13g2_decap_8
X_3451_ _0626_ _0624_ net609 _0627_ VPWR VGND sg13g2_mux2_1
X_3382_ _0550_ VPWR _0560_ VGND _0551_ _0559_ sg13g2_o21ai_1
X_5121_ _2060_ _2023_ _2059_ VPWR VGND sg13g2_xnor2_1
X_5052_ net724 net705 _1993_ VPWR VGND sg13g2_nor2_1
X_4003_ net1010 VPWR _1035_ VGND net883 _1021_ sg13g2_o21ai_1
XFILLER_19_891 VPWR VGND sg13g2_decap_8
X_4905_ _1849_ _1844_ _1848_ VPWR VGND sg13g2_nand2_1
X_4836_ _1404_ VPWR _1782_ VGND net1037 _1646_ sg13g2_o21ai_1
XFILLER_21_533 VPWR VGND sg13g2_decap_4
XFILLER_21_544 VPWR VGND sg13g2_decap_8
X_4767_ _1677_ _1713_ _1714_ VPWR VGND sg13g2_and2_1
X_3718_ _0877_ _0874_ _0875_ VPWR VGND sg13g2_nand2b_1
X_4698_ VPWR _1646_ _1645_ VGND sg13g2_inv_1
XFILLER_4_209 VPWR VGND sg13g2_fill_2
X_3649_ _0815_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] net608 VPWR VGND sg13g2_nand2_1
X_5319_ net63 VGND VPWR _0078_ ppwm_i.u_ppwm.pwm_value\[6\] clknet_leaf_16_clk sg13g2_dfrbpq_2
XFILLER_1_938 VPWR VGND sg13g2_decap_8
Xhold12 _0174_ VPWR VGND net384 sg13g2_dlygate4sd3_1
Xhold23 _0156_ VPWR VGND net395 sg13g2_dlygate4sd3_1
Xhold45 ppwm_i.u_ppwm.u_mem.memory\[82\] VPWR VGND net417 sg13g2_dlygate4sd3_1
Xhold34 _0283_ VPWR VGND net406 sg13g2_dlygate4sd3_1
Xhold56 falu_i.falutop.i2c_inst.op\[3\] VPWR VGND net428 sg13g2_dlygate4sd3_1
Xhold78 _0163_ VPWR VGND net450 sg13g2_dlygate4sd3_1
Xhold67 falu_i.falutop.div_inst.a\[6\] VPWR VGND net439 sg13g2_dlygate4sd3_1
XFILLER_21_1015 VPWR VGND sg13g2_decap_8
Xhold89 ppwm_i.u_ppwm.u_mem.memory\[109\] VPWR VGND net461 sg13g2_dlygate4sd3_1
XFILLER_28_121 VPWR VGND sg13g2_fill_1
XFILLER_44_603 VPWR VGND sg13g2_fill_1
XFILLER_28_165 VPWR VGND sg13g2_fill_2
XFILLER_43_113 VPWR VGND sg13g2_decap_4
XFILLER_43_102 VPWR VGND sg13g2_decap_8
XFILLER_25_883 VPWR VGND sg13g2_decap_8
XFILLER_12_555 VPWR VGND sg13g2_fill_2
XFILLER_40_875 VPWR VGND sg13g2_decap_8
XFILLER_8_515 VPWR VGND sg13g2_decap_8
X_5244__207 VPWR VGND net207 sg13g2_tiehi
XFILLER_0_960 VPWR VGND sg13g2_decap_8
XFILLER_48_942 VPWR VGND sg13g2_decap_8
XFILLER_47_474 VPWR VGND sg13g2_decap_8
XFILLER_19_198 VPWR VGND sg13g2_fill_2
X_2951_ _2305_ net750 VPWR VGND sg13g2_inv_2
XFILLER_43_691 VPWR VGND sg13g2_fill_2
X_2882_ _2236_ net1169 VPWR VGND sg13g2_inv_2
X_4621_ _1224_ _1507_ _1570_ VPWR VGND sg13g2_nor2_1
XFILLER_31_875 VPWR VGND sg13g2_fill_2
X_4552_ VGND VPWR _1363_ _1368_ _1502_ _1299_ sg13g2_a21oi_1
Xhold515 ppwm_i.u_ppwm.pwm_value\[9\] VPWR VGND net1167 sg13g2_dlygate4sd3_1
X_3503_ _0676_ VPWR _0677_ VGND _2246_ net597 sg13g2_o21ai_1
Xhold526 falu_i.falutop.data_in\[15\] VPWR VGND net1178 sg13g2_dlygate4sd3_1
X_4483_ _1379_ _1431_ _1433_ _1434_ VPWR VGND sg13g2_nor3_1
Xhold504 _1041_ VPWR VGND net1156 sg13g2_dlygate4sd3_1
X_3434_ net608 net611 _0610_ VPWR VGND sg13g2_nor2b_1
Xhold537 ppwm_i.u_ppwm.global_counter\[3\] VPWR VGND net1189 sg13g2_dlygate4sd3_1
X_3365_ _0543_ _0541_ _0542_ _2269_ ppwm_i.u_ppwm.pwm_value\[6\] VPWR VGND sg13g2_a22oi_1
X_3296_ _0478_ _2360_ VPWR VGND _2344_ sg13g2_nand2b_2
X_5104_ VGND VPWR _2305_ net564 _2044_ _1282_ sg13g2_a21oi_1
X_5035_ net815 VPWR _1977_ VGND net1020 net627 sg13g2_o21ai_1
XFILLER_26_669 VPWR VGND sg13g2_fill_2
XFILLER_15_36 VPWR VGND sg13g2_fill_2
XFILLER_22_831 VPWR VGND sg13g2_decap_8
X_4819_ _1763_ _1764_ _1758_ _1765_ VPWR VGND sg13g2_nand3_1
X_5386__280 VPWR VGND net280 sg13g2_tiehi
X_5527__165 VPWR VGND net165 sg13g2_tiehi
XFILLER_29_430 VPWR VGND sg13g2_decap_8
XFILLER_45_901 VPWR VGND sg13g2_decap_8
XFILLER_44_422 VPWR VGND sg13g2_fill_1
XFILLER_29_496 VPWR VGND sg13g2_decap_4
XFILLER_45_978 VPWR VGND sg13g2_decap_8
XFILLER_31_105 VPWR VGND sg13g2_decap_8
XFILLER_31_116 VPWR VGND sg13g2_fill_2
XFILLER_13_831 VPWR VGND sg13g2_decap_8
XFILLER_9_846 VPWR VGND sg13g2_decap_8
Xclkbuf_3_1__f_clk clknet_0_clk clknet_3_1__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_4_540 VPWR VGND sg13g2_decap_4
XFILLER_4_562 VPWR VGND sg13g2_decap_4
X_3150_ _2431_ _2439_ _0378_ VPWR VGND sg13g2_nor2_1
X_3081_ falu_i.falutop.i2c_inst.counter\[1\] falu_i.falutop.i2c_inst.counter\[0\]
+ _2432_ VPWR VGND sg13g2_and2_1
XFILLER_36_934 VPWR VGND sg13g2_decap_8
X_3983_ net808 VPWR _1020_ VGND net971 net652 sg13g2_o21ai_1
X_2934_ VPWR _2288_ net381 VGND sg13g2_inv_1
X_2865_ VPWR _2219_ net477 VGND sg13g2_inv_1
XFILLER_30_182 VPWR VGND sg13g2_fill_1
XFILLER_11_1014 VPWR VGND sg13g2_decap_8
X_4604_ _1485_ VPWR _1553_ VGND _1483_ _1486_ sg13g2_o21ai_1
Xhold301 _2095_ VPWR VGND net953 sg13g2_dlygate4sd3_1
X_2796_ VPWR _2150_ net411 VGND sg13g2_inv_1
X_5483__319 VPWR VGND net319 sg13g2_tiehi
X_4535_ net741 net762 net745 _1485_ VPWR VGND net756 sg13g2_nand4_1
Xhold334 _0349_ VPWR VGND net986 sg13g2_dlygate4sd3_1
Xhold312 falu_i.falutop.alu_inst.op\[3\] VPWR VGND net964 sg13g2_dlygate4sd3_1
Xhold323 _0448_ VPWR VGND net975 sg13g2_dlygate4sd3_1
Xhold356 ppwm_i.u_ppwm.u_mem.memory\[48\] VPWR VGND net1008 sg13g2_dlygate4sd3_1
Xhold378 _0310_ VPWR VGND net1030 sg13g2_dlygate4sd3_1
Xhold367 _0307_ VPWR VGND net1019 sg13g2_dlygate4sd3_1
X_4466_ _1416_ _1415_ _1417_ VPWR VGND sg13g2_nor2b_1
Xhold345 _1094_ VPWR VGND net997 sg13g2_dlygate4sd3_1
Xfanout825 net826 net825 VPWR VGND sg13g2_buf_8
X_3417_ VPWR VGND _2248_ _0594_ ppwm_i.u_ppwm.global_counter\[14\] _2247_ _0595_ ppwm_i.u_ppwm.global_counter\[15\]
+ sg13g2_a221oi_1
Xfanout803 net805 net803 VPWR VGND sg13g2_buf_8
Xhold389 falu_i.falutop.i2c_inst.result\[7\] VPWR VGND net1041 sg13g2_dlygate4sd3_1
X_4397_ VGND VPWR net628 _1348_ _0295_ _1349_ sg13g2_a21oi_1
Xfanout814 rst_n net814 VPWR VGND sg13g2_buf_8
X_3348_ VPWR VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] _0525_ _2247_ ppwm_i.u_ppwm.u_ex.reg_value_q\[6\]
+ _0526_ _2246_ sg13g2_a221oi_1
Xfanout836 net842 net836 VPWR VGND sg13g2_buf_8
X_3279_ _0462_ _2287_ ppwm_i.u_ppwm.u_pwm.counter\[1\] _2286_ ppwm_i.u_ppwm.u_pwm.counter\[2\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_38_282 VPWR VGND sg13g2_fill_2
X_5018_ _1960_ _1935_ _1959_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_945 VPWR VGND sg13g2_decap_8
XFILLER_14_617 VPWR VGND sg13g2_fill_2
XFILLER_14_639 VPWR VGND sg13g2_fill_2
XFILLER_42_959 VPWR VGND sg13g2_decap_8
XFILLER_10_845 VPWR VGND sg13g2_decap_8
XFILLER_21_160 VPWR VGND sg13g2_decap_4
XFILLER_22_683 VPWR VGND sg13g2_decap_4
XFILLER_5_348 VPWR VGND sg13g2_decap_8
XFILLER_1_521 VPWR VGND sg13g2_fill_2
XFILLER_29_260 VPWR VGND sg13g2_fill_1
XFILLER_18_956 VPWR VGND sg13g2_decap_8
XFILLER_45_797 VPWR VGND sg13g2_decap_4
XFILLER_17_488 VPWR VGND sg13g2_decap_8
XFILLER_32_425 VPWR VGND sg13g2_fill_2
XFILLER_32_447 VPWR VGND sg13g2_fill_1
XFILLER_16_90 VPWR VGND sg13g2_fill_2
XFILLER_34_1025 VPWR VGND sg13g2_decap_4
XFILLER_5_860 VPWR VGND sg13g2_decap_8
X_4320_ VGND VPWR _2296_ net750 _1273_ _1272_ sg13g2_a21oi_1
X_4251_ _1209_ net856 net607 VPWR VGND sg13g2_nand2_1
X_3202_ _0411_ net1060 net1090 VPWR VGND sg13g2_nand2_2
XFILLER_41_1018 VPWR VGND sg13g2_decap_8
X_4182_ _1157_ _1117_ _1118_ VPWR VGND sg13g2_xnor2_1
X_3133_ VGND VPWR net800 _0365_ _0014_ _0366_ sg13g2_a21oi_1
X_3064_ _2418_ _2414_ _2417_ _2410_ net786 VPWR VGND sg13g2_a22oi_1
XFILLER_35_285 VPWR VGND sg13g2_fill_1
XFILLER_35_296 VPWR VGND sg13g2_fill_2
X_3966_ VGND VPWR _2162_ net667 _0202_ _1011_ sg13g2_a21oi_1
X_2917_ _2271_ net1189 VPWR VGND sg13g2_inv_2
X_3897_ net840 VPWR _0977_ VGND net962 net649 sg13g2_o21ai_1
X_2848_ VPWR _2202_ net949 VGND sg13g2_inv_1
XFILLER_12_37 VPWR VGND sg13g2_fill_2
X_5567_ net89 VGND VPWR net1087 falu_i.falutop.alu_data_in\[13\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_2
XFILLER_3_819 VPWR VGND sg13g2_decap_8
Xhold120 ppwm_i.u_ppwm.u_pwm.cmp_value\[6\] VPWR VGND net492 sg13g2_dlygate4sd3_1
X_4518_ VGND VPWR net735 net721 _1468_ net760 sg13g2_a21oi_1
Xhold153 falu_i.falutop.div_inst.i\[0\] VPWR VGND net525 sg13g2_dlygate4sd3_1
X_5498_ net279 VGND VPWR _0257_ falu_i.falutop.div_inst.b1\[2\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
Xhold142 _0218_ VPWR VGND net514 sg13g2_dlygate4sd3_1
Xhold131 _0189_ VPWR VGND net503 sg13g2_dlygate4sd3_1
Xhold164 _0033_ VPWR VGND net536 sg13g2_dlygate4sd3_1
Xhold175 ppwm_i.u_ppwm.u_mem.memory\[33\] VPWR VGND net547 sg13g2_dlygate4sd3_1
Xhold186 _0157_ VPWR VGND net558 sg13g2_dlygate4sd3_1
X_4449_ VGND VPWR _1399_ _1400_ _1401_ _1362_ sg13g2_a21oi_1
Xfanout600 net604 net600 VPWR VGND sg13g2_buf_8
Xfanout611 net613 net611 VPWR VGND sg13g2_buf_8
Xfanout622 _1078_ net622 VPWR VGND sg13g2_buf_8
Xfanout633 net635 net633 VPWR VGND sg13g2_buf_8
Xhold197 _0228_ VPWR VGND net849 sg13g2_dlygate4sd3_1
Xfanout644 net645 net644 VPWR VGND sg13g2_buf_8
Xfanout666 net680 net666 VPWR VGND sg13g2_buf_8
Xfanout655 net666 net655 VPWR VGND sg13g2_buf_2
Xfanout677 net678 net677 VPWR VGND sg13g2_buf_8
Xfanout688 _2312_ net688 VPWR VGND sg13g2_buf_8
Xfanout699 _2309_ net699 VPWR VGND sg13g2_buf_8
XFILLER_2_1023 VPWR VGND sg13g2_decap_4
XFILLER_27_720 VPWR VGND sg13g2_decap_8
XFILLER_42_701 VPWR VGND sg13g2_fill_1
XFILLER_41_233 VPWR VGND sg13g2_fill_1
XFILLER_15_959 VPWR VGND sg13g2_decap_8
XFILLER_26_274 VPWR VGND sg13g2_decap_4
XFILLER_5_112 VPWR VGND sg13g2_fill_2
XFILLER_2_841 VPWR VGND sg13g2_decap_8
XFILLER_49_333 VPWR VGND sg13g2_decap_8
XFILLER_18_720 VPWR VGND sg13g2_fill_2
XFILLER_18_753 VPWR VGND sg13g2_fill_2
XFILLER_32_222 VPWR VGND sg13g2_fill_1
X_3820_ VGND VPWR _2214_ net643 _0129_ _0938_ sg13g2_a21oi_1
XFILLER_20_406 VPWR VGND sg13g2_decap_4
XFILLER_32_244 VPWR VGND sg13g2_fill_1
XFILLER_33_778 VPWR VGND sg13g2_decap_8
XFILLER_33_789 VPWR VGND sg13g2_decap_8
XFILLER_14_992 VPWR VGND sg13g2_decap_8
X_3751_ VGND VPWR _2293_ net686 _0094_ _0904_ sg13g2_a21oi_1
X_3682_ _0845_ _0702_ _0844_ VPWR VGND sg13g2_nand2_1
X_5421_ net208 VGND VPWR _0180_ ppwm_i.u_ppwm.u_mem.memory\[80\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_2
X_5352_ net348 VGND VPWR _0111_ ppwm_i.u_ppwm.u_mem.memory\[11\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_4303_ _1256_ _1222_ _1255_ VPWR VGND sg13g2_xnor2_1
X_5283_ net131 VGND VPWR _0045_ ppwm_i.u_ppwm.global_counter\[0\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_4234_ VGND VPWR net781 falu_i.falutop.div_inst.a\[4\] _1198_ _1197_ sg13g2_a21oi_1
X_4165_ VGND VPWR _2152_ net635 _0265_ net940 sg13g2_a21oi_1
X_3116_ VGND VPWR net802 _0353_ _0009_ _0354_ sg13g2_a21oi_1
X_4096_ net983 net999 net1054 net920 _1099_ VPWR VGND sg13g2_nor4_1
X_3047_ _2401_ net693 _2223_ net701 _2218_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_767 VPWR VGND sg13g2_decap_8
X_4998_ _1940_ _1937_ _1938_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_36 VPWR VGND sg13g2_decap_8
X_5489__303 VPWR VGND net303 sg13g2_tiehi
X_3949_ net840 VPWR _1003_ VGND net867 net674 sg13g2_o21ai_1
XFILLER_20_951 VPWR VGND sg13g2_decap_8
XFILLER_2_104 VPWR VGND sg13g2_fill_1
XFILLER_15_756 VPWR VGND sg13g2_fill_2
XFILLER_30_704 VPWR VGND sg13g2_fill_2
XFILLER_11_951 VPWR VGND sg13g2_decap_8
XFILLER_7_944 VPWR VGND sg13g2_decap_8
XFILLER_31_1017 VPWR VGND sg13g2_decap_8
XFILLER_31_1028 VPWR VGND sg13g2_fill_1
XFILLER_9_1007 VPWR VGND sg13g2_decap_8
XFILLER_49_141 VPWR VGND sg13g2_fill_2
X_4921_ _1856_ _1862_ _1864_ _1865_ VPWR VGND sg13g2_or3_1
X_4852_ _1797_ _1792_ _1796_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_704 VPWR VGND sg13g2_decap_8
XFILLER_21_726 VPWR VGND sg13g2_fill_1
X_3803_ net828 VPWR _0930_ VGND ppwm_i.u_ppwm.u_mem.memory\[21\] net661 sg13g2_o21ai_1
X_4783_ net720 net747 _1729_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_225 VPWR VGND sg13g2_fill_1
XFILLER_20_236 VPWR VGND sg13g2_fill_2
XFILLER_21_748 VPWR VGND sg13g2_decap_8
X_3734_ _0791_ net570 _0889_ _0891_ _0892_ VPWR VGND sg13g2_nor4_1
X_3665_ VPWR VGND _0656_ net799 _0829_ _2242_ _0083_ net570 sg13g2_a221oi_1
X_5404_ net244 VGND VPWR net450 ppwm_i.u_ppwm.u_mem.memory\[63\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_47_1002 VPWR VGND sg13g2_decap_8
X_3596_ _0765_ _2245_ net601 VPWR VGND sg13g2_xnor2_1
X_5335_ net33 VGND VPWR net468 falu_i.falutop.i2c_inst.op\[2\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_5266_ net164 VGND VPWR net471 ppwm_i.u_ppwm.u_pwm.cmp_value\[4\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
X_5345__362 VPWR VGND net362 sg13g2_tiehi
X_4217_ net779 _2152_ _1185_ VPWR VGND sg13g2_nor2_1
X_5197_ net777 VPWR _2114_ VGND falu_i.falutop.data_in\[0\] falu_i.falutop.data_in\[1\]
+ sg13g2_o21ai_1
X_4148_ net778 _1141_ net918 _0253_ VPWR VGND sg13g2_nor3_1
XFILLER_44_829 VPWR VGND sg13g2_fill_1
XFILLER_37_870 VPWR VGND sg13g2_fill_1
X_4079_ VPWR VGND falu_i.falutop.i2c_inst.result\[14\] _2154_ _0343_ falu_i.falutop.i2c_inst.result\[13\]
+ _1083_ _2445_ sg13g2_a221oi_1
XFILLER_28_358 VPWR VGND sg13g2_decap_8
XFILLER_43_339 VPWR VGND sg13g2_decap_8
XFILLER_34_13 VPWR VGND sg13g2_decap_8
XFILLER_11_203 VPWR VGND sg13g2_fill_2
XFILLER_34_57 VPWR VGND sg13g2_fill_2
XFILLER_12_759 VPWR VGND sg13g2_decap_4
Xclkload1 clknet_3_5__leaf_clk clkload1/X VPWR VGND sg13g2_buf_8
XFILLER_4_936 VPWR VGND sg13g2_decap_8
X_5396__260 VPWR VGND net260 sg13g2_tiehi
XFILLER_15_542 VPWR VGND sg13g2_fill_1
XFILLER_43_873 VPWR VGND sg13g2_fill_1
XFILLER_15_586 VPWR VGND sg13g2_decap_8
XFILLER_30_523 VPWR VGND sg13g2_fill_2
XFILLER_30_534 VPWR VGND sg13g2_fill_1
XFILLER_7_741 VPWR VGND sg13g2_decap_8
X_5548__285 VPWR VGND net285 sg13g2_tiehi
X_3450_ _0625_ VPWR _0626_ VGND _2249_ net595 sg13g2_o21ai_1
X_3381_ VPWR VGND _2239_ _0558_ ppwm_i.u_ppwm.global_counter\[4\] _2238_ _0559_ ppwm_i.u_ppwm.global_counter\[5\]
+ sg13g2_a221oi_1
XFILLER_3_980 VPWR VGND sg13g2_decap_8
X_5120_ VGND VPWR _2025_ _2026_ _2059_ _2058_ sg13g2_a21oi_1
X_5051_ _1803_ _1952_ _1992_ VPWR VGND sg13g2_nor2_1
XFILLER_38_612 VPWR VGND sg13g2_decap_4
X_4002_ _0215_ net808 _1033_ _1034_ VPWR VGND sg13g2_and3_1
XFILLER_38_678 VPWR VGND sg13g2_fill_2
XFILLER_19_870 VPWR VGND sg13g2_decap_8
X_4904_ _1848_ _1845_ _1846_ VPWR VGND sg13g2_xnor2_1
X_4835_ _1738_ _1780_ _1732_ _1781_ VPWR VGND sg13g2_nand3_1
X_4766_ _1711_ _1679_ _1712_ _1713_ VPWR VGND sg13g2_a21o_2
X_3717_ _0876_ _0875_ _0874_ VPWR VGND sg13g2_nand2b_1
X_4697_ net937 _1644_ _1645_ VPWR VGND sg13g2_nor2_1
X_3648_ _0814_ net419 VPWR VGND _0812_ sg13g2_nand2b_2
X_3579_ _0749_ _0747_ _0748_ VPWR VGND sg13g2_nand2_1
XFILLER_1_917 VPWR VGND sg13g2_decap_8
X_5318_ net65 VGND VPWR _0077_ ppwm_i.u_ppwm.pwm_value\[5\] clknet_leaf_13_clk sg13g2_dfrbpq_2
Xhold13 ppwm_i.u_ppwm.u_ex.state_q\[1\] VPWR VGND net385 sg13g2_dlygate4sd3_1
Xhold35 ppwm_i.u_ppwm.u_mem.memory\[50\] VPWR VGND net407 sg13g2_dlygate4sd3_1
Xhold46 _0181_ VPWR VGND net418 sg13g2_dlygate4sd3_1
Xhold24 falu_i.falutop.div_inst.acc_next\[0\] VPWR VGND net396 sg13g2_dlygate4sd3_1
X_5249_ net197 VGND VPWR _0011_ falu_i.falutop.i2c_inst.data_in\[7\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
XFILLER_29_57 VPWR VGND sg13g2_fill_2
Xhold68 _0342_ VPWR VGND net440 sg13g2_dlygate4sd3_1
Xhold57 _0095_ VPWR VGND net429 sg13g2_dlygate4sd3_1
XFILLER_28_111 VPWR VGND sg13g2_fill_1
Xhold79 ppwm_i.u_ppwm.u_mem.memory\[7\] VPWR VGND net451 sg13g2_dlygate4sd3_1
XFILLER_29_678 VPWR VGND sg13g2_fill_2
XFILLER_28_199 VPWR VGND sg13g2_decap_8
XFILLER_25_862 VPWR VGND sg13g2_decap_8
XFILLER_40_832 VPWR VGND sg13g2_fill_2
XFILLER_6_17 VPWR VGND sg13g2_fill_2
XFILLER_4_777 VPWR VGND sg13g2_fill_2
XFILLER_48_921 VPWR VGND sg13g2_decap_8
XFILLER_48_998 VPWR VGND sg13g2_decap_8
X_5578__289 VPWR VGND net289 sg13g2_tiehi
XFILLER_19_133 VPWR VGND sg13g2_decap_4
XFILLER_35_626 VPWR VGND sg13g2_fill_1
XFILLER_16_895 VPWR VGND sg13g2_decap_8
X_2950_ net766 _2304_ VPWR VGND sg13g2_inv_4
X_2881_ _2235_ net1160 VPWR VGND sg13g2_inv_2
XFILLER_31_854 VPWR VGND sg13g2_fill_1
X_4620_ _1568_ VPWR _1569_ VGND _1496_ _1566_ sg13g2_o21ai_1
X_4551_ _1288_ _1500_ net744 _1501_ VPWR VGND sg13g2_nand3_1
X_3502_ _0676_ ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] net596 VPWR VGND sg13g2_nand2_1
Xhold527 _0328_ VPWR VGND net1179 sg13g2_dlygate4sd3_1
X_4482_ VGND VPWR net737 net769 _1433_ _1430_ sg13g2_a21oi_1
Xhold505 _0217_ VPWR VGND net1157 sg13g2_dlygate4sd3_1
Xhold516 ppwm_i.u_ppwm.pc\[1\] VPWR VGND net1168 sg13g2_dlygate4sd3_1
Xhold538 ppwm_i.u_ppwm.pwm_value\[7\] VPWR VGND net1190 sg13g2_dlygate4sd3_1
X_3433_ net598 net608 _0609_ VPWR VGND sg13g2_nor2_1
X_3364_ _0542_ ppwm_i.u_ppwm.global_counter\[5\] _2247_ ppwm_i.u_ppwm.global_counter\[6\]
+ _2246_ VPWR VGND sg13g2_a22oi_1
X_5103_ _2040_ _2041_ _1317_ _2043_ VPWR VGND _2042_ sg13g2_nand4_1
X_3295_ _0477_ _2257_ net599 VPWR VGND sg13g2_xnor2_1
X_5034_ net627 _1975_ _1976_ VPWR VGND sg13g2_and2_1
XFILLER_39_987 VPWR VGND sg13g2_decap_8
XFILLER_38_497 VPWR VGND sg13g2_fill_2
XFILLER_41_607 VPWR VGND sg13g2_decap_8
XFILLER_40_106 VPWR VGND sg13g2_decap_8
XFILLER_22_810 VPWR VGND sg13g2_decap_8
XFILLER_22_887 VPWR VGND sg13g2_decap_8
X_4818_ _1759_ VPWR _1764_ VGND _1760_ _1762_ sg13g2_o21ai_1
X_4749_ _1696_ net757 net733 net762 net728 VPWR VGND sg13g2_a22oi_1
XFILLER_0_202 VPWR VGND sg13g2_decap_4
XFILLER_1_714 VPWR VGND sg13g2_fill_1
XFILLER_1_725 VPWR VGND sg13g2_fill_2
XFILLER_49_718 VPWR VGND sg13g2_decap_8
XFILLER_5_1021 VPWR VGND sg13g2_decap_8
XFILLER_29_453 VPWR VGND sg13g2_decap_4
XFILLER_44_401 VPWR VGND sg13g2_fill_1
XFILLER_17_615 VPWR VGND sg13g2_fill_1
XFILLER_29_475 VPWR VGND sg13g2_decap_8
XFILLER_45_957 VPWR VGND sg13g2_decap_8
XFILLER_16_147 VPWR VGND sg13g2_fill_2
XFILLER_13_887 VPWR VGND sg13g2_decap_8
XFILLER_4_552 VPWR VGND sg13g2_fill_1
X_3080_ _2431_ net1016 _2430_ VPWR VGND sg13g2_nand2_2
X_5402__248 VPWR VGND net248 sg13g2_tiehi
X_3982_ VGND VPWR _2156_ net668 _0210_ _1019_ sg13g2_a21oi_1
X_2933_ VPWR _2287_ net506 VGND sg13g2_inv_1
X_2864_ VPWR _2218_ net402 VGND sg13g2_inv_1
X_5583_ net231 VGND VPWR net440 falu_i.falutop.div_inst.a\[6\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_2795_ VPWR _2149_ net435 VGND sg13g2_inv_1
X_4603_ _1549_ _1551_ _1552_ VPWR VGND sg13g2_nor2_1
X_4534_ net745 net741 net763 net757 _1484_ VPWR VGND sg13g2_and4_1
Xhold302 ppwm_i.u_ppwm.global_counter\[11\] VPWR VGND net954 sg13g2_dlygate4sd3_1
Xhold324 _0059_ VPWR VGND net976 sg13g2_dlygate4sd3_1
Xhold335 _0350_ VPWR VGND net987 sg13g2_dlygate4sd3_1
Xhold313 ppwm_i.u_ppwm.u_mem.memory\[21\] VPWR VGND net965 sg13g2_dlygate4sd3_1
Xhold357 falu_i.falutop.div_inst.acc\[0\] VPWR VGND net1009 sg13g2_dlygate4sd3_1
Xhold368 falu_i.falutop.i2c_inst.result\[11\] VPWR VGND net1020 sg13g2_dlygate4sd3_1
X_4465_ VGND VPWR net735 net725 _1416_ net765 sg13g2_a21oi_1
Xhold346 _0244_ VPWR VGND net998 sg13g2_dlygate4sd3_1
Xhold379 ppwm_i.u_ppwm.global_counter\[19\] VPWR VGND net1031 sg13g2_dlygate4sd3_1
X_3416_ VPWR VGND ppwm_i.u_ppwm.pwm_value\[3\] _0593_ _2264_ ppwm_i.u_ppwm.pwm_value\[4\]
+ _0594_ _2263_ sg13g2_a221oi_1
Xfanout815 net817 net815 VPWR VGND sg13g2_buf_8
X_4396_ net818 VPWR _1349_ VGND net1022 net628 sg13g2_o21ai_1
Xfanout804 net805 net804 VPWR VGND sg13g2_buf_8
X_3347_ VPWR VGND _2239_ _0524_ ppwm_i.u_ppwm.pwm_value\[4\] _2238_ _0525_ ppwm_i.u_ppwm.pwm_value\[5\]
+ sg13g2_a221oi_1
Xfanout837 net838 net837 VPWR VGND sg13g2_buf_8
Xfanout826 net832 net826 VPWR VGND sg13g2_buf_2
X_5017_ _1957_ _1943_ _1959_ VPWR VGND sg13g2_xor2_1
X_3278_ _0460_ VPWR _0461_ VGND ppwm_i.u_ppwm.u_pwm.counter\[0\] _2288_ sg13g2_o21ai_1
XFILLER_38_261 VPWR VGND sg13g2_decap_8
XFILLER_26_14 VPWR VGND sg13g2_fill_2
XFILLER_27_924 VPWR VGND sg13g2_decap_8
XFILLER_38_294 VPWR VGND sg13g2_decap_4
XFILLER_26_25 VPWR VGND sg13g2_fill_2
XFILLER_42_938 VPWR VGND sg13g2_decap_8
XFILLER_13_139 VPWR VGND sg13g2_decap_8
XFILLER_21_183 VPWR VGND sg13g2_fill_1
XFILLER_1_500 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_27_1022 VPWR VGND sg13g2_decap_8
XFILLER_18_935 VPWR VGND sg13g2_decap_8
XFILLER_44_231 VPWR VGND sg13g2_decap_4
XFILLER_45_787 VPWR VGND sg13g2_fill_1
XFILLER_44_264 VPWR VGND sg13g2_fill_2
XFILLER_17_456 VPWR VGND sg13g2_decap_4
XFILLER_34_1004 VPWR VGND sg13g2_decap_8
XFILLER_13_695 VPWR VGND sg13g2_decap_8
XFILLER_9_655 VPWR VGND sg13g2_decap_8
X_5285__127 VPWR VGND net127 sg13g2_tiehi
XFILLER_4_393 VPWR VGND sg13g2_fill_1
XFILLER_4_371 VPWR VGND sg13g2_fill_1
X_4250_ _1208_ VPWR _0289_ VGND _1098_ _1163_ sg13g2_o21ai_1
X_4181_ VGND VPWR net634 _1155_ _0272_ _1156_ sg13g2_a21oi_1
X_3201_ VGND VPWR _2277_ _0407_ _0038_ _0410_ sg13g2_a21oi_1
X_3132_ net816 VPWR _0366_ VGND net945 _0365_ sg13g2_o21ai_1
XFILLER_27_209 VPWR VGND sg13g2_fill_1
X_3063_ VGND VPWR _2415_ _2416_ _2417_ net786 sg13g2_a21oi_1
XFILLER_36_732 VPWR VGND sg13g2_decap_4
XFILLER_24_949 VPWR VGND sg13g2_decap_8
X_3965_ net836 VPWR _1011_ VGND ppwm_i.u_ppwm.u_mem.memory\[102\] net667 sg13g2_o21ai_1
X_3896_ VGND VPWR _2187_ net678 _0167_ _0976_ sg13g2_a21oi_1
XFILLER_32_982 VPWR VGND sg13g2_decap_8
X_2916_ _2270_ net1107 VPWR VGND sg13g2_inv_2
X_2847_ VPWR _2201_ net434 VGND sg13g2_inv_1
Xhold110 ppwm_i.u_ppwm.u_mem.memory\[72\] VPWR VGND net482 sg13g2_dlygate4sd3_1
X_5566_ net100 VGND VPWR net1104 falu_i.falutop.alu_data_in\[12\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_2
Xhold121 _0030_ VPWR VGND net493 sg13g2_dlygate4sd3_1
X_4517_ net735 net760 _1467_ VPWR VGND sg13g2_and2_1
X_5497_ net281 VGND VPWR _0256_ falu_i.falutop.div_inst.b1\[1\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
Xhold143 ppwm_i.u_ppwm.u_mem.memory\[16\] VPWR VGND net515 sg13g2_dlygate4sd3_1
Xhold132 ppwm_i.u_ppwm.u_mem.memory\[10\] VPWR VGND net504 sg13g2_dlygate4sd3_1
Xhold176 _0133_ VPWR VGND net548 sg13g2_dlygate4sd3_1
Xhold154 _1139_ VPWR VGND net526 sg13g2_dlygate4sd3_1
X_4448_ VGND VPWR _1308_ _1398_ _1400_ _1310_ sg13g2_a21oi_1
Xhold165 ppwm_i.u_ppwm.u_mem.memory\[99\] VPWR VGND net537 sg13g2_dlygate4sd3_1
Xfanout601 net604 net601 VPWR VGND sg13g2_buf_8
Xfanout612 net613 net612 VPWR VGND sg13g2_buf_1
Xfanout623 net624 net623 VPWR VGND sg13g2_buf_8
Xhold198 falu_i.falutop.i2c_inst.data_in\[6\] VPWR VGND net850 sg13g2_dlygate4sd3_1
Xhold187 ppwm_i.u_ppwm.u_mem.memory\[110\] VPWR VGND net559 sg13g2_dlygate4sd3_1
Xfanout656 net658 net656 VPWR VGND sg13g2_buf_8
Xfanout645 net651 net645 VPWR VGND sg13g2_buf_8
Xfanout634 net635 net634 VPWR VGND sg13g2_buf_8
X_4379_ net743 net740 _1332_ VPWR VGND sg13g2_nor2_1
Xfanout667 net668 net667 VPWR VGND sg13g2_buf_8
Xfanout678 net679 net678 VPWR VGND sg13g2_buf_8
Xfanout689 _2312_ net689 VPWR VGND sg13g2_buf_1
XFILLER_2_1002 VPWR VGND sg13g2_decap_8
XFILLER_41_201 VPWR VGND sg13g2_fill_2
XFILLER_15_938 VPWR VGND sg13g2_decap_8
X_5355__342 VPWR VGND net342 sg13g2_tiehi
XFILLER_41_267 VPWR VGND sg13g2_decap_8
XFILLER_23_982 VPWR VGND sg13g2_decap_8
XFILLER_10_632 VPWR VGND sg13g2_decap_4
XFILLER_6_614 VPWR VGND sg13g2_fill_1
XFILLER_5_102 VPWR VGND sg13g2_fill_1
XFILLER_2_820 VPWR VGND sg13g2_decap_8
XFILLER_2_897 VPWR VGND sg13g2_decap_8
XFILLER_17_231 VPWR VGND sg13g2_fill_2
XFILLER_33_735 VPWR VGND sg13g2_fill_2
XFILLER_32_234 VPWR VGND sg13g2_fill_1
XFILLER_14_971 VPWR VGND sg13g2_decap_8
X_3750_ falu_i.falutop.i2c_inst.data_in\[18\] net686 _0904_ VPWR VGND sg13g2_nor2_1
XFILLER_32_267 VPWR VGND sg13g2_decap_8
XFILLER_9_441 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_fill_1
XFILLER_13_481 VPWR VGND sg13g2_fill_1
X_3681_ VGND VPWR net577 _0843_ _0844_ net569 sg13g2_a21oi_1
X_5420_ net212 VGND VPWR _0179_ ppwm_i.u_ppwm.u_mem.memory\[79\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_5351_ net350 VGND VPWR _0110_ ppwm_i.u_ppwm.u_mem.memory\[10\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
XFILLER_5_691 VPWR VGND sg13g2_fill_2
X_4302_ _1253_ _1225_ _1255_ VPWR VGND sg13g2_xor2_1
X_5282_ net132 VGND VPWR net865 ppwm_i.u_ppwm.period_start clknet_leaf_12_clk sg13g2_dfrbpq_2
X_4233_ net781 _2148_ _1197_ VPWR VGND sg13g2_nor2_1
X_4164_ net803 VPWR _1147_ VGND net939 net635 sg13g2_o21ai_1
X_4095_ _1098_ _1095_ VPWR VGND _1096_ sg13g2_nand2b_2
X_3115_ net804 VPWR _0354_ VGND net869 _0353_ sg13g2_o21ai_1
X_3046_ VPWR VGND _2204_ _2399_ net693 _2213_ _2400_ net699 sg13g2_a221oi_1
XFILLER_23_201 VPWR VGND sg13g2_decap_8
XFILLER_24_746 VPWR VGND sg13g2_decap_8
X_4997_ net727 net706 _1937_ _1939_ VPWR VGND sg13g2_nor3_1
XFILLER_23_15 VPWR VGND sg13g2_decap_8
XFILLER_23_289 VPWR VGND sg13g2_decap_8
XFILLER_20_930 VPWR VGND sg13g2_decap_8
XFILLER_32_790 VPWR VGND sg13g2_decap_8
X_3948_ VGND VPWR _2169_ net672 _0193_ _1002_ sg13g2_a21oi_1
X_3879_ net839 VPWR _0968_ VGND net866 net676 sg13g2_o21ai_1
XFILLER_3_617 VPWR VGND sg13g2_decap_8
X_5549_ net259 VGND VPWR net1036 falu_i.falutop.i2c_inst.result\[13\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_3_639 VPWR VGND sg13g2_decap_8
XFILLER_15_713 VPWR VGND sg13g2_decap_4
XFILLER_27_584 VPWR VGND sg13g2_decap_8
XFILLER_14_223 VPWR VGND sg13g2_fill_2
X_5472__341 VPWR VGND net341 sg13g2_tiehi
XFILLER_42_587 VPWR VGND sg13g2_fill_1
XFILLER_11_930 VPWR VGND sg13g2_decap_8
XFILLER_7_923 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_4
X_5307__87 VPWR VGND net87 sg13g2_tiehi
X_5322__57 VPWR VGND net57 sg13g2_tiehi
XFILLER_36_7 VPWR VGND sg13g2_fill_2
X_4920_ VGND VPWR _1860_ _1861_ _1864_ _1857_ sg13g2_a21oi_1
XFILLER_18_595 VPWR VGND sg13g2_decap_4
X_4851_ _1796_ _1653_ _1793_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_738 VPWR VGND sg13g2_fill_2
X_3802_ VGND VPWR _2220_ net653 _0120_ _0929_ sg13g2_a21oi_1
X_4782_ VGND VPWR _1242_ _1726_ _1728_ _1727_ sg13g2_a21oi_1
X_3733_ VGND VPWR net582 _0794_ _0891_ _0890_ sg13g2_a21oi_1
X_3664_ _0665_ net570 _0826_ _0828_ _0829_ VPWR VGND sg13g2_nor4_1
X_5403_ net246 VGND VPWR _0162_ ppwm_i.u_ppwm.u_mem.memory\[62\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_3595_ VPWR VGND _0764_ net798 _0752_ _2246_ _0078_ net572 sg13g2_a221oi_1
X_5334_ net34 VGND VPWR net913 falu_i.falutop.i2c_inst.op\[1\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_2
X_5265_ net166 VGND VPWR net458 ppwm_i.u_ppwm.u_pwm.cmp_value\[3\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_1
X_4216_ VGND VPWR net634 _1183_ _0279_ net1080 sg13g2_a21oi_1
X_5196_ net891 net624 _2113_ VPWR VGND sg13g2_nor2_1
X_4147_ net917 _1138_ _1142_ VPWR VGND sg13g2_nor2_1
X_4078_ _1082_ _2438_ falu_i.falutop.i2c_inst.result\[12\] _2432_ falu_i.falutop.i2c_inst.result\[15\]
+ VPWR VGND sg13g2_a22oi_1
X_3029_ VGND VPWR _2207_ net688 _2383_ net708 sg13g2_a21oi_1
XFILLER_24_532 VPWR VGND sg13g2_fill_2
XFILLER_34_47 VPWR VGND sg13g2_fill_1
XFILLER_11_237 VPWR VGND sg13g2_decap_8
XFILLER_12_749 VPWR VGND sg13g2_fill_2
Xclkload2 clknet_3_7__leaf_clk clkload2/X VPWR VGND sg13g2_buf_8
XFILLER_4_915 VPWR VGND sg13g2_decap_8
XFILLER_46_123 VPWR VGND sg13g2_fill_1
XFILLER_43_830 VPWR VGND sg13g2_fill_2
XFILLER_28_871 VPWR VGND sg13g2_decap_8
XFILLER_43_841 VPWR VGND sg13g2_fill_2
XFILLER_42_340 VPWR VGND sg13g2_fill_2
XFILLER_42_384 VPWR VGND sg13g2_fill_1
XFILLER_24_91 VPWR VGND sg13g2_fill_2
XFILLER_30_579 VPWR VGND sg13g2_decap_4
XFILLER_6_241 VPWR VGND sg13g2_decap_4
X_3380_ _0558_ _0552_ _0557_ _2270_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_34_4 VPWR VGND sg13g2_decap_4
XFILLER_2_491 VPWR VGND sg13g2_fill_1
X_5050_ _1991_ _1988_ _1989_ VPWR VGND sg13g2_xnor2_1
X_4001_ _1034_ net1186 _1030_ VPWR VGND sg13g2_nand2_1
X_4903_ _1847_ _1846_ _1845_ VPWR VGND sg13g2_nand2b_1
XFILLER_18_381 VPWR VGND sg13g2_fill_2
XFILLER_33_373 VPWR VGND sg13g2_decap_8
X_4834_ _1780_ _1779_ net615 _1725_ _1723_ VPWR VGND sg13g2_a22oi_1
X_5412__228 VPWR VGND net228 sg13g2_tiehi
XFILLER_14_1013 VPWR VGND sg13g2_decap_8
X_4765_ net615 VPWR _1712_ VGND _1679_ _1711_ sg13g2_o21ai_1
XFILLER_21_557 VPWR VGND sg13g2_fill_2
XFILLER_21_568 VPWR VGND sg13g2_decap_8
X_3716_ VGND VPWR ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] net601 _0875_ _0868_ sg13g2_a21oi_1
X_4696_ _1585_ _1404_ _1644_ VPWR VGND sg13g2_nor2b_1
X_3647_ _2255_ _0812_ _0813_ VPWR VGND sg13g2_nor2_2
X_3578_ _0748_ _0712_ _0729_ VPWR VGND sg13g2_nand2_1
X_5317_ net67 VGND VPWR net1182 ppwm_i.u_ppwm.pwm_value\[4\] clknet_leaf_18_clk sg13g2_dfrbpq_2
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_0_439 VPWR VGND sg13g2_decap_8
Xhold14 _2426_ VPWR VGND net386 sg13g2_dlygate4sd3_1
Xhold36 _0150_ VPWR VGND net408 sg13g2_dlygate4sd3_1
Xhold47 ppwm_i.u_ppwm.u_ex.state_q\[2\] VPWR VGND net419 sg13g2_dlygate4sd3_1
Xhold25 _0286_ VPWR VGND net397 sg13g2_dlygate4sd3_1
X_5248_ net199 VGND VPWR _0010_ falu_i.falutop.i2c_inst.data_in\[6\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
Xhold58 ppwm_i.u_ppwm.u_pwm.cmp_value\[7\] VPWR VGND net430 sg13g2_dlygate4sd3_1
X_5179_ VGND VPWR net705 net619 _0320_ _2106_ sg13g2_a21oi_1
XFILLER_29_624 VPWR VGND sg13g2_fill_2
Xhold69 ppwm_i.u_ppwm.u_mem.memory\[8\] VPWR VGND net441 sg13g2_dlygate4sd3_1
XFILLER_40_800 VPWR VGND sg13g2_fill_1
XFILLER_4_734 VPWR VGND sg13g2_decap_8
XFILLER_3_255 VPWR VGND sg13g2_fill_1
XFILLER_48_900 VPWR VGND sg13g2_decap_8
XFILLER_0_995 VPWR VGND sg13g2_decap_8
XFILLER_48_977 VPWR VGND sg13g2_decap_8
XFILLER_19_80 VPWR VGND sg13g2_fill_1
XFILLER_37_1013 VPWR VGND sg13g2_decap_8
XFILLER_16_874 VPWR VGND sg13g2_decap_8
XFILLER_15_384 VPWR VGND sg13g2_fill_2
X_2880_ VPWR _2234_ net523 VGND sg13g2_inv_1
XFILLER_42_192 VPWR VGND sg13g2_fill_1
XFILLER_31_877 VPWR VGND sg13g2_fill_1
X_4550_ _1295_ _1298_ _1500_ VPWR VGND sg13g2_nor2_1
Xhold517 ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] VPWR VGND net1169 sg13g2_dlygate4sd3_1
XFILLER_7_594 VPWR VGND sg13g2_decap_8
Xhold506 falu_i.falutop.data_in\[8\] VPWR VGND net1158 sg13g2_dlygate4sd3_1
X_4481_ VPWR _1432_ _1431_ VGND sg13g2_inv_1
X_3501_ net602 net574 _0674_ _0675_ VPWR VGND sg13g2_nor3_1
Xhold539 _0079_ VPWR VGND net1191 sg13g2_dlygate4sd3_1
X_3432_ _2345_ _2360_ _0608_ VPWR VGND sg13g2_and2_1
Xhold528 ppwm_i.u_ppwm.global_counter\[15\] VPWR VGND net1180 sg13g2_dlygate4sd3_1
X_3363_ _0540_ VPWR _0541_ VGND _2247_ ppwm_i.u_ppwm.global_counter\[5\] sg13g2_o21ai_1
XFILLER_44_1028 VPWR VGND sg13g2_fill_1
X_5102_ _2042_ _2005_ _2039_ VPWR VGND sg13g2_nand2_1
X_3294_ _0476_ net793 net599 VPWR VGND sg13g2_nand2_1
XFILLER_38_421 VPWR VGND sg13g2_fill_1
X_5033_ _1973_ _1974_ net638 _1975_ VPWR VGND sg13g2_nand3_1
XFILLER_39_966 VPWR VGND sg13g2_decap_8
X_5295__107 VPWR VGND net107 sg13g2_tiehi
X_5452__78 VPWR VGND net78 sg13g2_tiehi
X_4817_ _1759_ _1760_ _1762_ _1763_ VPWR VGND sg13g2_or3_1
XFILLER_22_866 VPWR VGND sg13g2_decap_8
X_4748_ net728 net762 net732 _1695_ VPWR VGND net756 sg13g2_nand4_1
XFILLER_31_37 VPWR VGND sg13g2_fill_2
X_4679_ _1627_ _1626_ VPWR VGND _1625_ sg13g2_nand2b_2
XFILLER_0_225 VPWR VGND sg13g2_fill_1
XFILLER_5_1000 VPWR VGND sg13g2_decap_8
XFILLER_45_936 VPWR VGND sg13g2_decap_8
XFILLER_44_457 VPWR VGND sg13g2_decap_8
XFILLER_12_343 VPWR VGND sg13g2_fill_2
XFILLER_13_866 VPWR VGND sg13g2_decap_8
X_5365__322 VPWR VGND net322 sg13g2_tiehi
XFILLER_39_229 VPWR VGND sg13g2_fill_2
XFILLER_0_792 VPWR VGND sg13g2_decap_8
XFILLER_35_402 VPWR VGND sg13g2_fill_2
XFILLER_36_969 VPWR VGND sg13g2_decap_8
X_3981_ net836 VPWR _1019_ VGND net559 net668 sg13g2_o21ai_1
X_2932_ VPWR _2286_ net520 VGND sg13g2_inv_1
Xclkbuf_leaf_42_clk clknet_3_1__leaf_clk clknet_leaf_42_clk VPWR VGND sg13g2_buf_8
XFILLER_15_181 VPWR VGND sg13g2_fill_1
X_2863_ VPWR _2217_ net950 VGND sg13g2_inv_1
X_5582_ net239 VGND VPWR net466 falu_i.falutop.div_inst.a\[5\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_2794_ VPWR _2148_ net405 VGND sg13g2_inv_1
X_4602_ _1551_ net752 net745 net770 net728 VPWR VGND sg13g2_a22oi_1
XFILLER_8_881 VPWR VGND sg13g2_decap_8
X_4533_ _1483_ net737 net767 VPWR VGND sg13g2_nand2_1
Xhold325 ppwm_i.u_ppwm.u_mem.memory\[73\] VPWR VGND net977 sg13g2_dlygate4sd3_1
XFILLER_7_94 VPWR VGND sg13g2_fill_2
Xhold303 _0443_ VPWR VGND net955 sg13g2_dlygate4sd3_1
Xhold314 _0120_ VPWR VGND net966 sg13g2_dlygate4sd3_1
Xhold369 _0306_ VPWR VGND net1021 sg13g2_dlygate4sd3_1
X_4464_ net725 net765 net735 _1415_ VPWR VGND sg13g2_nand3_1
Xhold347 falu_i.falutop.div_inst.b\[4\] VPWR VGND net999 sg13g2_dlygate4sd3_1
Xhold336 _0351_ VPWR VGND net988 sg13g2_dlygate4sd3_1
Xhold358 ppwm_i.u_ppwm.u_mem.bit_count\[4\] VPWR VGND net1010 sg13g2_dlygate4sd3_1
X_4395_ _1347_ VPWR _1348_ VGND falu_i.falutop.div_inst.val\[0\] _1074_ sg13g2_o21ai_1
Xfanout805 net806 net805 VPWR VGND sg13g2_buf_8
Xfanout816 net817 net816 VPWR VGND sg13g2_buf_8
X_3415_ VPWR VGND _2250_ _0592_ ppwm_i.u_ppwm.global_counter\[12\] _2249_ _0593_ ppwm_i.u_ppwm.global_counter\[13\]
+ sg13g2_a221oi_1
Xfanout838 net841 net838 VPWR VGND sg13g2_buf_8
Xfanout827 net831 net827 VPWR VGND sg13g2_buf_8
X_3346_ VPWR VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] _0523_ _2249_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\]
+ _0524_ _2248_ sg13g2_a221oi_1
X_5016_ _1943_ _1957_ _1958_ VPWR VGND sg13g2_nor2_1
XFILLER_27_903 VPWR VGND sg13g2_decap_8
X_3277_ _0460_ ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] ppwm_i.u_ppwm.u_pwm.counter\[1\]
+ VPWR VGND sg13g2_nand2b_1
XFILLER_38_284 VPWR VGND sg13g2_fill_1
XFILLER_14_619 VPWR VGND sg13g2_fill_1
XFILLER_41_449 VPWR VGND sg13g2_fill_1
XFILLER_41_427 VPWR VGND sg13g2_decap_4
XFILLER_35_991 VPWR VGND sg13g2_decap_8
XFILLER_22_652 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_33_clk clknet_3_6__leaf_clk clknet_leaf_33_clk VPWR VGND sg13g2_buf_8
XFILLER_21_151 VPWR VGND sg13g2_decap_4
XFILLER_27_1001 VPWR VGND sg13g2_decap_8
XFILLER_49_516 VPWR VGND sg13g2_fill_2
XFILLER_45_711 VPWR VGND sg13g2_fill_1
XFILLER_18_914 VPWR VGND sg13g2_decap_8
XFILLER_29_240 VPWR VGND sg13g2_fill_2
XFILLER_44_221 VPWR VGND sg13g2_decap_4
XFILLER_33_939 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_24_clk clknet_3_6__leaf_clk clknet_leaf_24_clk VPWR VGND sg13g2_buf_8
XFILLER_9_601 VPWR VGND sg13g2_fill_1
XFILLER_13_652 VPWR VGND sg13g2_fill_2
XFILLER_25_490 VPWR VGND sg13g2_fill_2
XFILLER_41_983 VPWR VGND sg13g2_decap_8
XFILLER_9_678 VPWR VGND sg13g2_decap_8
X_5482__321 VPWR VGND net321 sg13g2_tiehi
XFILLER_5_895 VPWR VGND sg13g2_decap_8
X_3200_ _0410_ net809 _0409_ VPWR VGND sg13g2_nand2_1
X_4180_ net803 VPWR _1156_ VGND net1116 net634 sg13g2_o21ai_1
X_3131_ _0344_ _0360_ _0365_ VPWR VGND sg13g2_nor2_1
X_3062_ VPWR VGND _2227_ net790 net688 _2232_ _2416_ net696 sg13g2_a221oi_1
XFILLER_36_700 VPWR VGND sg13g2_fill_1
XFILLER_24_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_15_clk clknet_3_2__leaf_clk clknet_leaf_15_clk VPWR VGND sg13g2_buf_8
X_3964_ VGND VPWR _2163_ net668 _0201_ _1010_ sg13g2_a21oi_1
XFILLER_32_961 VPWR VGND sg13g2_decap_8
X_3895_ net839 VPWR _0976_ VGND net889 net676 sg13g2_o21ai_1
X_2915_ _2269_ net1184 VPWR VGND sg13g2_inv_2
X_2846_ _2200_ net407 VPWR VGND sg13g2_inv_2
XFILLER_12_39 VPWR VGND sg13g2_fill_1
Xhold100 ppwm_i.u_ppwm.u_mem.memory\[35\] VPWR VGND net472 sg13g2_dlygate4sd3_1
X_5565_ net108 VGND VPWR net1102 falu_i.falutop.alu_data_in\[11\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_2
Xhold144 ppwm_i.u_ppwm.u_mem.memory\[31\] VPWR VGND net516 sg13g2_dlygate4sd3_1
X_4516_ _1466_ net740 net716 VPWR VGND sg13g2_nand2_1
Xhold122 falu_i.falutop.div_inst.acc\[3\] VPWR VGND net494 sg13g2_dlygate4sd3_1
X_5496_ net283 VGND VPWR _0255_ falu_i.falutop.div_inst.b1\[0\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
Xhold111 ppwm_i.u_ppwm.u_mem.memory\[6\] VPWR VGND net483 sg13g2_dlygate4sd3_1
Xhold133 _0109_ VPWR VGND net505 sg13g2_dlygate4sd3_1
Xhold177 falu_i.falutop.div_inst.acc\[5\] VPWR VGND net549 sg13g2_dlygate4sd3_1
Xhold155 _0252_ VPWR VGND net527 sg13g2_dlygate4sd3_1
X_4447_ VGND VPWR _1399_ _1398_ _1308_ sg13g2_or2_1
Xhold166 _0199_ VPWR VGND net538 sg13g2_dlygate4sd3_1
Xfanout602 net604 net602 VPWR VGND sg13g2_buf_8
Xfanout613 _2389_ net613 VPWR VGND sg13g2_buf_1
Xfanout624 net626 net624 VPWR VGND sg13g2_buf_1
Xhold199 _0234_ VPWR VGND net851 sg13g2_dlygate4sd3_1
Xhold188 ppwm_i.u_ppwm.u_mem.memory\[4\] VPWR VGND net560 sg13g2_dlygate4sd3_1
Xfanout657 net658 net657 VPWR VGND sg13g2_buf_1
Xfanout635 _1134_ net635 VPWR VGND sg13g2_buf_8
X_4378_ VGND VPWR net707 _1330_ _1331_ net743 sg13g2_a21oi_1
Xfanout646 net651 net646 VPWR VGND sg13g2_buf_8
X_3329_ _2373_ _0507_ _0508_ VPWR VGND sg13g2_nor2_1
Xfanout679 net680 net679 VPWR VGND sg13g2_buf_8
Xfanout668 net679 net668 VPWR VGND sg13g2_buf_2
XFILLER_39_582 VPWR VGND sg13g2_fill_2
XFILLER_15_917 VPWR VGND sg13g2_decap_8
XFILLER_41_213 VPWR VGND sg13g2_fill_1
XFILLER_14_416 VPWR VGND sg13g2_decap_8
XFILLER_23_961 VPWR VGND sg13g2_decap_8
XFILLER_10_600 VPWR VGND sg13g2_decap_4
X_5319__63 VPWR VGND net63 sg13g2_tiehi
XFILLER_6_648 VPWR VGND sg13g2_decap_4
XFILLER_10_688 VPWR VGND sg13g2_fill_1
XFILLER_2_876 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_decap_8
XFILLER_27_80 VPWR VGND sg13g2_fill_1
XFILLER_32_202 VPWR VGND sg13g2_fill_1
XFILLER_14_950 VPWR VGND sg13g2_decap_8
X_3680_ ppwm_i.u_ppwm.pwm_value\[3\] _0704_ net581 _0843_ VPWR VGND sg13g2_mux2_1
XFILLER_9_497 VPWR VGND sg13g2_decap_8
X_5350_ net352 VGND VPWR net505 ppwm_i.u_ppwm.u_mem.memory\[9\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_5281_ net134 VGND VPWR net1025 ppwm_i.u_ppwm.u_pwm.counter\[9\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
XFILLER_5_670 VPWR VGND sg13g2_fill_2
X_4301_ _1225_ _1253_ _1254_ VPWR VGND sg13g2_and2_1
XFILLER_4_40 VPWR VGND sg13g2_fill_1
X_4232_ VGND VPWR _1106_ _1195_ _0283_ _1196_ sg13g2_a21oi_1
Xclkbuf_leaf_4_clk clknet_3_3__leaf_clk clknet_leaf_4_clk VPWR VGND sg13g2_buf_8
X_4163_ _1145_ _1146_ _0264_ VPWR VGND sg13g2_nor2_1
X_4094_ _1096_ _1095_ _1097_ VPWR VGND sg13g2_nor2b_2
X_3114_ _2446_ net987 _0353_ VPWR VGND sg13g2_nor2_1
XFILLER_49_880 VPWR VGND sg13g2_decap_8
X_3045_ ppwm_i.u_ppwm.u_mem.memory\[38\] _2313_ _2399_ VPWR VGND sg13g2_nor2_1
X_5519__206 VPWR VGND net206 sg13g2_tiehi
XFILLER_24_725 VPWR VGND sg13g2_decap_8
X_4996_ net727 net705 _1938_ VPWR VGND sg13g2_nor2_1
XFILLER_12_909 VPWR VGND sg13g2_decap_8
XFILLER_11_419 VPWR VGND sg13g2_fill_2
X_3947_ net838 VPWR _1002_ VGND net401 net672 sg13g2_o21ai_1
X_3878_ VGND VPWR _2194_ net670 _0158_ _0967_ sg13g2_a21oi_1
XFILLER_20_986 VPWR VGND sg13g2_decap_8
X_2829_ VPWR _2183_ net922 VGND sg13g2_inv_1
X_5548_ net285 VGND VPWR net1019 falu_i.falutop.i2c_inst.result\[12\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_5479_ net327 VGND VPWR net946 falu_i.falutop.data_in\[10\] clknet_leaf_7_clk sg13g2_dfrbpq_2
XFILLER_24_1026 VPWR VGND sg13g2_fill_2
XFILLER_47_817 VPWR VGND sg13g2_fill_2
XFILLER_46_338 VPWR VGND sg13g2_fill_1
XFILLER_7_902 VPWR VGND sg13g2_decap_8
XFILLER_6_401 VPWR VGND sg13g2_fill_1
XFILLER_11_986 VPWR VGND sg13g2_decap_8
XFILLER_13_60 VPWR VGND sg13g2_fill_1
XFILLER_7_979 VPWR VGND sg13g2_decap_8
X_5251__193 VPWR VGND net193 sg13g2_tiehi
XFILLER_2_651 VPWR VGND sg13g2_decap_8
XFILLER_49_198 VPWR VGND sg13g2_decap_8
XFILLER_18_541 VPWR VGND sg13g2_decap_8
XFILLER_18_552 VPWR VGND sg13g2_fill_1
Xclkbuf_3_7__f_clk clknet_0_clk clknet_3_7__leaf_clk VPWR VGND sg13g2_buf_8
X_4850_ VPWR _1795_ _1794_ VGND sg13g2_inv_1
X_3801_ net827 VPWR _0929_ VGND ppwm_i.u_ppwm.u_mem.memory\[20\] net653 sg13g2_o21ai_1
X_4781_ _1373_ VPWR _1727_ VGND net632 _1726_ sg13g2_o21ai_1
XFILLER_20_238 VPWR VGND sg13g2_fill_1
X_3732_ net580 VPWR _0890_ VGND ppwm_i.u_ppwm.pwm_value\[8\] net583 sg13g2_o21ai_1
X_3663_ VGND VPWR net582 _0662_ _0828_ _0827_ sg13g2_a21oi_1
X_5402_ net248 VGND VPWR _0161_ ppwm_i.u_ppwm.u_mem.memory\[61\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_3594_ net572 _0759_ _0763_ _0764_ VPWR VGND sg13g2_nor3_1
XFILLER_6_990 VPWR VGND sg13g2_decap_8
X_5333_ net35 VGND VPWR net421 falu_i.falutop.i2c_inst.op\[0\] clknet_leaf_7_clk sg13g2_dfrbpq_1
X_5264_ net168 VGND VPWR net521 ppwm_i.u_ppwm.u_pwm.cmp_value\[2\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
X_4215_ net805 VPWR _1184_ VGND net1079 net635 sg13g2_o21ai_1
X_5195_ _2110_ VPWR _0330_ VGND net622 _2112_ sg13g2_o21ai_1
X_4146_ net409 _1140_ _1141_ VPWR VGND sg13g2_nor2_1
XFILLER_28_316 VPWR VGND sg13g2_decap_8
X_4077_ VPWR VGND falu_i.falutop.i2c_inst.result\[8\] _1079_ _2438_ falu_i.falutop.i2c_inst.result\[11\]
+ _1081_ _2432_ sg13g2_a221oi_1
X_3028_ ppwm_i.u_ppwm.u_mem.memory\[33\] net791 net793 _2382_ VPWR VGND sg13g2_nor3_1
XFILLER_37_883 VPWR VGND sg13g2_fill_1
XFILLER_11_205 VPWR VGND sg13g2_fill_1
XFILLER_24_566 VPWR VGND sg13g2_fill_2
XFILLER_34_59 VPWR VGND sg13g2_fill_1
X_4979_ _1922_ _1878_ _1880_ _1920_ VPWR VGND sg13g2_and3_1
XFILLER_12_739 VPWR VGND sg13g2_decap_4
Xclkload3 VPWR clkload3/Y clknet_leaf_44_clk VGND sg13g2_inv_1
XFILLER_20_783 VPWR VGND sg13g2_fill_1
XFILLER_19_327 VPWR VGND sg13g2_fill_2
XFILLER_15_533 VPWR VGND sg13g2_decap_8
XFILLER_15_555 VPWR VGND sg13g2_fill_1
XFILLER_7_776 VPWR VGND sg13g2_decap_4
XFILLER_7_754 VPWR VGND sg13g2_fill_2
XFILLER_7_787 VPWR VGND sg13g2_fill_1
X_5543__36 VPWR VGND net36 sg13g2_tiehi
X_5509__249 VPWR VGND net249 sg13g2_tiehi
X_4000_ _1033_ _1032_ _1030_ VPWR VGND sg13g2_nand2b_1
XFILLER_38_658 VPWR VGND sg13g2_fill_1
XFILLER_26_809 VPWR VGND sg13g2_decap_8
X_5375__302 VPWR VGND net302 sg13g2_tiehi
XFILLER_34_820 VPWR VGND sg13g2_decap_8
X_4902_ net738 net706 _1846_ VPWR VGND sg13g2_nor2_1
XFILLER_33_341 VPWR VGND sg13g2_fill_1
X_4833_ _1778_ _1739_ _1779_ VPWR VGND sg13g2_xor2_1
X_4764_ _1709_ _1680_ _1711_ VPWR VGND sg13g2_xor2_1
X_3715_ _0874_ _2236_ net601 VPWR VGND sg13g2_xnor2_1
X_4695_ _1642_ VPWR _1643_ VGND _1604_ _1606_ sg13g2_o21ai_1
X_3646_ _0812_ _0811_ net579 _0612_ net598 VPWR VGND sg13g2_a22oi_1
X_3577_ net600 VPWR _0747_ VGND ppwm_i.u_ppwm.pwm_value\[5\] ppwm_i.u_ppwm.pwm_value\[4\]
+ sg13g2_o21ai_1
XFILLER_0_418 VPWR VGND sg13g2_decap_8
X_5316_ net69 VGND VPWR _0075_ ppwm_i.u_ppwm.pwm_value\[3\] clknet_leaf_12_clk sg13g2_dfrbpq_2
X_5247_ net201 VGND VPWR _0009_ falu_i.falutop.i2c_inst.data_in\[5\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
Xhold26 ppwm_i.u_ppwm.u_mem.memory\[55\] VPWR VGND net398 sg13g2_dlygate4sd3_1
Xhold37 falu_i.falutop.div_inst.i\[2\] VPWR VGND net409 sg13g2_dlygate4sd3_1
Xhold15 _0001_ VPWR VGND net387 sg13g2_dlygate4sd3_1
Xhold59 _0031_ VPWR VGND net431 sg13g2_dlygate4sd3_1
X_5178_ net1137 net619 _2106_ VPWR VGND sg13g2_nor2_1
Xhold48 falu_i.falutop.i2c_inst.op\[0\] VPWR VGND net420 sg13g2_dlygate4sd3_1
X_4129_ net879 _1130_ _1131_ VPWR VGND sg13g2_nor2_1
XFILLER_29_658 VPWR VGND sg13g2_fill_2
XFILLER_12_536 VPWR VGND sg13g2_decap_8
XFILLER_24_385 VPWR VGND sg13g2_decap_8
XFILLER_25_897 VPWR VGND sg13g2_decap_8
XFILLER_12_547 VPWR VGND sg13g2_fill_2
XFILLER_8_529 VPWR VGND sg13g2_decap_4
XFILLER_6_19 VPWR VGND sg13g2_fill_1
XFILLER_4_779 VPWR VGND sg13g2_fill_1
XFILLER_10_50 VPWR VGND sg13g2_fill_2
XFILLER_3_289 VPWR VGND sg13g2_decap_8
XFILLER_0_974 VPWR VGND sg13g2_decap_8
XFILLER_19_113 VPWR VGND sg13g2_fill_2
XFILLER_48_956 VPWR VGND sg13g2_decap_8
XFILLER_47_444 VPWR VGND sg13g2_decap_8
XFILLER_47_433 VPWR VGND sg13g2_decap_8
XFILLER_19_146 VPWR VGND sg13g2_decap_8
XFILLER_16_853 VPWR VGND sg13g2_decap_8
X_3500_ _0673_ VPWR _0674_ VGND net584 _0630_ sg13g2_o21ai_1
Xhold518 _0089_ VPWR VGND net1170 sg13g2_dlygate4sd3_1
Xhold507 _0321_ VPWR VGND net1159 sg13g2_dlygate4sd3_1
X_4480_ _1431_ net737 net769 _1430_ VPWR VGND sg13g2_and3_2
X_3431_ VGND VPWR _2252_ _0606_ _0071_ _0607_ sg13g2_a21oi_1
Xhold529 ppwm_i.u_ppwm.pwm_value\[4\] VPWR VGND net1181 sg13g2_dlygate4sd3_1
X_3362_ VGND VPWR ppwm_i.u_ppwm.pwm_value\[4\] _2270_ _0540_ _0539_ sg13g2_a21oi_1
XFILLER_44_1007 VPWR VGND sg13g2_decap_8
X_5101_ _2041_ _2009_ _2039_ VPWR VGND sg13g2_nand2_1
X_3293_ VGND VPWR net376 _0474_ _0065_ _0475_ sg13g2_a21oi_1
X_5032_ falu_i.falutop.div_inst.rem\[3\] _1929_ net773 _1974_ VPWR VGND sg13g2_nand3_1
XFILLER_22_845 VPWR VGND sg13g2_decap_8
XFILLER_34_672 VPWR VGND sg13g2_decap_4
XFILLER_34_694 VPWR VGND sg13g2_decap_8
X_4816_ VGND VPWR net728 net758 _1762_ falu_i.falutop.alu_data_in\[7\] sg13g2_a21oi_1
XFILLER_33_193 VPWR VGND sg13g2_decap_8
X_4747_ net732 net728 net762 net756 _1694_ VPWR VGND sg13g2_and4_1
X_4678_ _1621_ VPWR _1626_ VGND _1623_ _1624_ sg13g2_o21ai_1
X_3629_ net573 _0791_ _0796_ _0797_ VPWR VGND sg13g2_nor3_1
XFILLER_1_727 VPWR VGND sg13g2_fill_1
XFILLER_29_411 VPWR VGND sg13g2_decap_8
XFILLER_45_915 VPWR VGND sg13g2_decap_8
XFILLER_16_105 VPWR VGND sg13g2_decap_4
XFILLER_17_606 VPWR VGND sg13g2_fill_2
XFILLER_17_628 VPWR VGND sg13g2_decap_8
XFILLER_17_639 VPWR VGND sg13g2_fill_1
XFILLER_13_801 VPWR VGND sg13g2_decap_8
XFILLER_25_672 VPWR VGND sg13g2_fill_1
XFILLER_40_631 VPWR VGND sg13g2_fill_1
XFILLER_13_845 VPWR VGND sg13g2_decap_8
X_5469__347 VPWR VGND net347 sg13g2_tiehi
XFILLER_4_532 VPWR VGND sg13g2_fill_2
XFILLER_47_230 VPWR VGND sg13g2_fill_2
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_36_948 VPWR VGND sg13g2_decap_8
XFILLER_23_609 VPWR VGND sg13g2_decap_8
X_3980_ VGND VPWR _2157_ net667 _0209_ _1018_ sg13g2_a21oi_1
X_2931_ VPWR _2285_ net457 VGND sg13g2_inv_1
Xclkbuf_0_clk clk clknet_0_clk VPWR VGND sg13g2_buf_8
X_4601_ VPWR _1550_ _1549_ VGND sg13g2_inv_1
XFILLER_30_163 VPWR VGND sg13g2_fill_1
X_2862_ VPWR _2216_ net508 VGND sg13g2_inv_1
X_2793_ VPWR _2147_ net432 VGND sg13g2_inv_1
X_5581_ net247 VGND VPWR net453 falu_i.falutop.div_inst.a\[4\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_8_860 VPWR VGND sg13g2_decap_8
XFILLER_11_1028 VPWR VGND sg13g2_fill_1
X_4532_ _1482_ net732 net769 VPWR VGND sg13g2_nand2_1
XFILLER_7_392 VPWR VGND sg13g2_decap_4
Xhold326 falu_i.falutop.div_inst.val\[2\] VPWR VGND net978 sg13g2_dlygate4sd3_1
X_4463_ _1414_ net743 net716 VPWR VGND sg13g2_nand2_1
Xhold315 falu_i.falutop.div_inst.b\[3\] VPWR VGND net967 sg13g2_dlygate4sd3_1
Xhold304 _0056_ VPWR VGND net956 sg13g2_dlygate4sd3_1
Xhold337 ppwm_i.u_ppwm.global_counter\[17\] VPWR VGND net989 sg13g2_dlygate4sd3_1
Xhold348 _0333_ VPWR VGND net1000 sg13g2_dlygate4sd3_1
Xhold359 _1035_ VPWR VGND net1011 sg13g2_dlygate4sd3_1
X_3414_ VPWR VGND net784 _0591_ _2266_ ppwm_i.u_ppwm.pwm_value\[2\] _0592_ _2265_
+ sg13g2_a221oi_1
X_4394_ _1347_ _1262_ _1346_ VPWR VGND sg13g2_nand2_1
Xfanout806 net814 net806 VPWR VGND sg13g2_buf_8
Xfanout839 net840 net839 VPWR VGND sg13g2_buf_8
Xfanout817 net823 net817 VPWR VGND sg13g2_buf_8
Xfanout828 net831 net828 VPWR VGND sg13g2_buf_2
X_3345_ VPWR VGND _2241_ _0522_ ppwm_i.u_ppwm.pwm_value\[2\] _2240_ _0523_ ppwm_i.u_ppwm.pwm_value\[3\]
+ sg13g2_a221oi_1
X_3276_ VGND VPWR _2258_ _0457_ _0064_ _0459_ sg13g2_a21oi_1
XFILLER_39_731 VPWR VGND sg13g2_fill_2
X_5015_ _1955_ _1946_ _1957_ VPWR VGND sg13g2_xor2_1
XFILLER_38_241 VPWR VGND sg13g2_decap_4
XFILLER_26_27 VPWR VGND sg13g2_fill_1
XFILLER_27_959 VPWR VGND sg13g2_decap_8
XFILLER_35_970 VPWR VGND sg13g2_decap_8
XFILLER_10_804 VPWR VGND sg13g2_decap_4
XFILLER_10_859 VPWR VGND sg13g2_decap_8
X_5401__250 VPWR VGND net250 sg13g2_tiehi
XFILLER_29_274 VPWR VGND sg13g2_decap_8
XFILLER_29_296 VPWR VGND sg13g2_decap_8
XFILLER_41_962 VPWR VGND sg13g2_decap_8
XFILLER_40_461 VPWR VGND sg13g2_decap_8
XFILLER_13_675 VPWR VGND sg13g2_decap_4
X_5337__31 VPWR VGND net31 sg13g2_tiehi
XFILLER_5_874 VPWR VGND sg13g2_decap_8
X_3130_ VGND VPWR net800 _0363_ _0013_ _0364_ sg13g2_a21oi_1
X_5261__173 VPWR VGND net173 sg13g2_tiehi
X_3061_ _2415_ net692 _2222_ net700 _2217_ VPWR VGND sg13g2_a22oi_1
XFILLER_35_222 VPWR VGND sg13g2_decap_4
XFILLER_24_907 VPWR VGND sg13g2_decap_8
XFILLER_17_981 VPWR VGND sg13g2_decap_8
X_3963_ net836 VPWR _1010_ VGND net500 net667 sg13g2_o21ai_1
XFILLER_32_940 VPWR VGND sg13g2_decap_8
X_3894_ VGND VPWR _2188_ net676 _0166_ _0975_ sg13g2_a21oi_1
X_2914_ _2268_ net1092 VPWR VGND sg13g2_inv_2
X_2845_ VPWR _2199_ net915 VGND sg13g2_inv_1
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_31_494 VPWR VGND sg13g2_fill_2
XFILLER_12_29 VPWR VGND sg13g2_fill_1
X_5564_ net116 VGND VPWR _0323_ falu_i.falutop.alu_data_in\[10\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
Xhold101 _0135_ VPWR VGND net473 sg13g2_dlygate4sd3_1
X_4515_ _1415_ VPWR _1465_ VGND _1416_ _1418_ sg13g2_o21ai_1
X_5495_ net287 VGND VPWR net410 falu_i.falutop.div_inst.i\[2\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
Xhold123 _0289_ VPWR VGND net495 sg13g2_dlygate4sd3_1
Xhold134 ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] VPWR VGND net506 sg13g2_dlygate4sd3_1
Xhold112 _0105_ VPWR VGND net484 sg13g2_dlygate4sd3_1
Xhold145 _0130_ VPWR VGND net517 sg13g2_dlygate4sd3_1
X_4446_ _1398_ _1395_ _1396_ VPWR VGND sg13g2_xnor2_1
Xhold167 ppwm_i.u_ppwm.u_mem.memory\[102\] VPWR VGND net539 sg13g2_dlygate4sd3_1
Xhold156 ppwm_i.u_ppwm.u_mem.memory\[106\] VPWR VGND net528 sg13g2_dlygate4sd3_1
Xfanout603 net604 net603 VPWR VGND sg13g2_buf_2
X_5383__286 VPWR VGND net286 sg13g2_tiehi
Xfanout614 _1590_ net614 VPWR VGND sg13g2_buf_8
Xhold178 _0291_ VPWR VGND net550 sg13g2_dlygate4sd3_1
X_4377_ _1330_ net730 net736 VPWR VGND sg13g2_nand2b_1
Xhold189 _0103_ VPWR VGND net561 sg13g2_dlygate4sd3_1
Xfanout658 net666 net658 VPWR VGND sg13g2_buf_8
Xfanout647 net651 net647 VPWR VGND sg13g2_buf_1
Xfanout625 net626 net625 VPWR VGND sg13g2_buf_8
Xfanout636 net637 net636 VPWR VGND sg13g2_buf_8
X_3328_ _2254_ _2367_ _0507_ VPWR VGND sg13g2_nor2_1
Xfanout669 net670 net669 VPWR VGND sg13g2_buf_8
X_3259_ VGND VPWR ppwm_i.u_ppwm.global_counter\[13\] _0445_ _0448_ net974 sg13g2_a21oi_1
XFILLER_27_734 VPWR VGND sg13g2_decap_4
XFILLER_26_233 VPWR VGND sg13g2_fill_1
XFILLER_41_203 VPWR VGND sg13g2_fill_1
XFILLER_23_940 VPWR VGND sg13g2_decap_8
XFILLER_10_656 VPWR VGND sg13g2_fill_2
X_5334__34 VPWR VGND net34 sg13g2_tiehi
XFILLER_2_855 VPWR VGND sg13g2_decap_8
XFILLER_1_321 VPWR VGND sg13g2_fill_1
XFILLER_1_354 VPWR VGND sg13g2_fill_1
XFILLER_49_358 VPWR VGND sg13g2_decap_8
XFILLER_33_704 VPWR VGND sg13g2_fill_2
XFILLER_33_715 VPWR VGND sg13g2_decap_8
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_13_494 VPWR VGND sg13g2_decap_8
X_5280_ net136 VGND VPWR net1095 ppwm_i.u_ppwm.u_pwm.counter\[8\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_2
XFILLER_5_693 VPWR VGND sg13g2_fill_1
X_4300_ _1253_ _1230_ _1252_ VPWR VGND sg13g2_xnor2_1
X_4231_ net405 net605 _1196_ VPWR VGND sg13g2_nor2_1
X_5523__182 VPWR VGND net182 sg13g2_tiehi
X_4162_ net803 VPWR _1146_ VGND net1133 net634 sg13g2_o21ai_1
X_4093_ _1096_ falu_i.falutop.div_inst.busy VPWR VGND net778 sg13g2_nand2b_2
X_3113_ VGND VPWR net800 net988 _0008_ _0352_ sg13g2_a21oi_1
X_3044_ VGND VPWR _2199_ net704 _2398_ net708 sg13g2_a21oi_1
XFILLER_24_704 VPWR VGND sg13g2_decap_8
XFILLER_36_531 VPWR VGND sg13g2_fill_1
XFILLER_36_564 VPWR VGND sg13g2_fill_2
X_4995_ _1937_ net723 net748 VPWR VGND sg13g2_nand2_1
XFILLER_17_1023 VPWR VGND sg13g2_decap_4
X_3946_ VGND VPWR _2170_ net648 _0192_ _1001_ sg13g2_a21oi_1
X_3877_ net834 VPWR _0967_ VGND net557 net670 sg13g2_o21ai_1
XFILLER_20_965 VPWR VGND sg13g2_decap_8
X_2828_ _2182_ net383 VPWR VGND sg13g2_inv_2
X_5547_ net293 VGND VPWR net1021 falu_i.falutop.i2c_inst.result\[11\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_2_118 VPWR VGND sg13g2_decap_8
X_5478_ net329 VGND VPWR net900 falu_i.falutop.data_in\[9\] clknet_leaf_37_clk sg13g2_dfrbpq_2
X_5465__361 VPWR VGND net361 sg13g2_tiehi
X_4429_ _1318_ _1378_ _1380_ _1381_ VPWR VGND sg13g2_nor3_1
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_24_1005 VPWR VGND sg13g2_decap_8
XFILLER_47_829 VPWR VGND sg13g2_fill_1
XFILLER_15_704 VPWR VGND sg13g2_fill_2
XFILLER_42_545 VPWR VGND sg13g2_decap_4
XFILLER_11_965 VPWR VGND sg13g2_decap_8
XFILLER_7_958 VPWR VGND sg13g2_decap_8
XFILLER_10_497 VPWR VGND sg13g2_decap_4
XFILLER_2_685 VPWR VGND sg13g2_fill_1
XFILLER_36_9 VPWR VGND sg13g2_fill_1
XFILLER_49_111 VPWR VGND sg13g2_decap_8
XFILLER_37_317 VPWR VGND sg13g2_decap_4
XFILLER_18_520 VPWR VGND sg13g2_decap_8
XFILLER_46_851 VPWR VGND sg13g2_fill_1
XFILLER_46_895 VPWR VGND sg13g2_decap_8
XFILLER_33_512 VPWR VGND sg13g2_decap_8
XFILLER_33_523 VPWR VGND sg13g2_fill_1
X_4780_ VGND VPWR _1246_ _1669_ _1726_ _1243_ sg13g2_a21oi_1
X_3800_ VGND VPWR _2221_ net641 _0119_ _0928_ sg13g2_a21oi_1
X_3731_ _0888_ _0887_ _0889_ VPWR VGND sg13g2_nor2b_1
XFILLER_9_251 VPWR VGND sg13g2_decap_8
X_3662_ net579 VPWR _0827_ VGND net785 net582 sg13g2_o21ai_1
X_5401_ net250 VGND VPWR net438 ppwm_i.u_ppwm.u_mem.memory\[60\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_3593_ VGND VPWR net588 _0761_ _0763_ _0762_ sg13g2_a21oi_1
X_5332_ net37 VGND VPWR net1161 ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_2
XFILLER_47_1027 VPWR VGND sg13g2_fill_2
XFILLER_47_1016 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_5263_ net170 VGND VPWR net507 ppwm_i.u_ppwm.u_pwm.cmp_value\[1\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_1
X_4214_ VPWR _1183_ _1182_ VGND sg13g2_inv_1
X_5194_ _2111_ falu_i.falutop.data_in\[1\] _2112_ VPWR VGND sg13g2_xor2_1
X_4145_ _1140_ net917 _1138_ VPWR VGND sg13g2_nand2_1
XFILLER_18_17 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_fill_2
X_4076_ VGND VPWR falu_i.falutop.i2c_inst.result\[9\] _2445_ _1080_ falu_i.falutop.i2c_inst.counter\[2\]
+ sg13g2_a21oi_1
XFILLER_43_309 VPWR VGND sg13g2_decap_4
X_3027_ VPWR VGND _2380_ _2254_ _2379_ _2376_ _2381_ _2378_ sg13g2_a221oi_1
X_4978_ VGND VPWR _1878_ _1880_ _1921_ _1920_ sg13g2_a21oi_1
XFILLER_20_751 VPWR VGND sg13g2_decap_8
X_3929_ net837 VPWR _0993_ VGND net878 net673 sg13g2_o21ai_1
Xclkload4 clkload4/Y clknet_leaf_18_clk VPWR VGND sg13g2_inv_8
XFILLER_3_449 VPWR VGND sg13g2_fill_2
XFILLER_3_438 VPWR VGND sg13g2_decap_8
XFILLER_8_1021 VPWR VGND sg13g2_decap_8
XFILLER_34_309 VPWR VGND sg13g2_decap_8
XFILLER_42_342 VPWR VGND sg13g2_fill_1
XFILLER_11_740 VPWR VGND sg13g2_decap_4
XFILLER_11_784 VPWR VGND sg13g2_decap_8
XFILLER_40_92 VPWR VGND sg13g2_decap_8
XFILLER_41_7 VPWR VGND sg13g2_decap_8
XFILLER_3_994 VPWR VGND sg13g2_decap_8
X_5479__327 VPWR VGND net327 sg13g2_tiehi
XFILLER_38_637 VPWR VGND sg13g2_decap_4
XFILLER_1_64 VPWR VGND sg13g2_fill_1
X_5555__215 VPWR VGND net215 sg13g2_tiehi
X_5950_ ppwm_i.u_ppwm.data_o net7 VPWR VGND sg13g2_buf_2
XFILLER_19_884 VPWR VGND sg13g2_decap_8
X_4901_ _1845_ net733 net748 VPWR VGND sg13g2_nand2_1
X_4832_ _1776_ _1708_ _1778_ VPWR VGND sg13g2_xor2_1
XFILLER_21_526 VPWR VGND sg13g2_decap_8
XFILLER_21_537 VPWR VGND sg13g2_fill_2
X_4763_ _1680_ _1709_ _1710_ VPWR VGND sg13g2_nor2_1
X_3714_ VPWR VGND _0873_ net798 _0870_ _2237_ _0088_ net569 sg13g2_a221oi_1
X_4694_ VPWR VGND net615 _1619_ _1641_ net616 _1642_ _1608_ sg13g2_a221oi_1
X_3645_ net612 _0609_ _0811_ VPWR VGND sg13g2_nor2_1
X_3576_ _0746_ _2246_ net601 VPWR VGND sg13g2_xnor2_1
X_5315_ net71 VGND VPWR _0074_ ppwm_i.u_ppwm.pwm_value\[2\] clknet_leaf_9_clk sg13g2_dfrbpq_2
X_5246_ net203 VGND VPWR _0008_ falu_i.falutop.i2c_inst.data_in\[4\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
Xhold38 _0254_ VPWR VGND net410 sg13g2_dlygate4sd3_1
Xhold27 falu_i.falutop.div_inst.quo\[1\] VPWR VGND net399 sg13g2_dlygate4sd3_1
Xhold16 falu_i.falutop.div_inst.a\[1\] VPWR VGND net388 sg13g2_dlygate4sd3_1
X_5177_ net1073 net749 net618 _0319_ VPWR VGND sg13g2_mux2_1
XFILLER_21_1008 VPWR VGND sg13g2_decap_8
Xhold49 _0092_ VPWR VGND net421 sg13g2_dlygate4sd3_1
X_4128_ _1110_ _1129_ _1130_ VPWR VGND sg13g2_nor2_1
XFILLER_45_15 VPWR VGND sg13g2_fill_1
X_5455__66 VPWR VGND net66 sg13g2_tiehi
X_4059_ net848 falu_i.falutop.data_in\[0\] net684 _0228_ VPWR VGND sg13g2_mux2_1
XFILLER_43_117 VPWR VGND sg13g2_fill_2
XFILLER_24_342 VPWR VGND sg13g2_fill_2
XFILLER_25_876 VPWR VGND sg13g2_decap_8
XFILLER_36_191 VPWR VGND sg13g2_decap_8
XFILLER_20_570 VPWR VGND sg13g2_decap_8
XFILLER_4_769 VPWR VGND sg13g2_decap_4
XFILLER_0_953 VPWR VGND sg13g2_decap_8
XFILLER_48_935 VPWR VGND sg13g2_decap_8
XFILLER_47_467 VPWR VGND sg13g2_decap_8
XFILLER_16_832 VPWR VGND sg13g2_decap_8
XFILLER_43_684 VPWR VGND sg13g2_decap_8
XFILLER_31_868 VPWR VGND sg13g2_decap_8
X_5411__230 VPWR VGND net230 sg13g2_tiehi
XFILLER_30_356 VPWR VGND sg13g2_fill_2
Xhold508 ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] VPWR VGND net1160 sg13g2_dlygate4sd3_1
X_3430_ net813 VPWR _0607_ VGND net592 _0606_ sg13g2_o21ai_1
Xhold519 ppwm_i.u_ppwm.pwm_value\[2\] VPWR VGND net1171 sg13g2_dlygate4sd3_1
X_3361_ VPWR VGND _2249_ _0538_ ppwm_i.u_ppwm.global_counter\[3\] _2248_ _0539_ ppwm_i.u_ppwm.global_counter\[4\]
+ sg13g2_a221oi_1
XFILLER_3_780 VPWR VGND sg13g2_fill_1
X_5100_ _2005_ _2009_ _2039_ _2040_ VPWR VGND sg13g2_or3_1
X_3292_ net810 VPWR _0475_ VGND net376 _0474_ sg13g2_o21ai_1
X_5031_ _1929_ net773 falu_i.falutop.div_inst.rem\[3\] _1973_ VPWR VGND sg13g2_a21o_1
X_5342__368 VPWR VGND net368 sg13g2_tiehi
XFILLER_38_445 VPWR VGND sg13g2_decap_4
XFILLER_22_824 VPWR VGND sg13g2_decap_8
X_4815_ falu_i.falutop.alu_data_in\[7\] net755 net727 _1761_ VPWR VGND sg13g2_nand3_1
X_4746_ _1693_ net723 net767 VPWR VGND sg13g2_nand2_1
X_4677_ _1621_ _1623_ _1624_ _1625_ VPWR VGND sg13g2_nor3_1
X_3628_ VGND VPWR net589 _0794_ _0796_ _0795_ sg13g2_a21oi_1
X_3559_ _0708_ _0712_ _0729_ _0730_ VPWR VGND sg13g2_or3_1
X_5229_ net452 net625 _2137_ VPWR VGND sg13g2_nor2_1
XFILLER_29_489 VPWR VGND sg13g2_decap_8
XFILLER_44_415 VPWR VGND sg13g2_decap_8
X_5393__266 VPWR VGND net266 sg13g2_tiehi
XFILLER_13_824 VPWR VGND sg13g2_decap_8
XFILLER_24_150 VPWR VGND sg13g2_decap_4
XFILLER_12_345 VPWR VGND sg13g2_fill_1
XFILLER_24_183 VPWR VGND sg13g2_fill_2
XFILLER_24_194 VPWR VGND sg13g2_decap_8
XFILLER_9_839 VPWR VGND sg13g2_decap_8
XFILLER_21_83 VPWR VGND sg13g2_decap_4
XFILLER_0_750 VPWR VGND sg13g2_decap_8
X_5248__199 VPWR VGND net199 sg13g2_tiehi
XFILLER_48_721 VPWR VGND sg13g2_fill_2
XFILLER_35_415 VPWR VGND sg13g2_decap_4
XFILLER_44_993 VPWR VGND sg13g2_decap_8
X_2930_ VPWR _2284_ net470 VGND sg13g2_inv_1
XFILLER_16_673 VPWR VGND sg13g2_decap_4
XFILLER_16_695 VPWR VGND sg13g2_fill_2
XFILLER_22_109 VPWR VGND sg13g2_fill_2
XFILLER_30_120 VPWR VGND sg13g2_decap_4
X_2861_ VPWR _2215_ net959 VGND sg13g2_inv_1
X_4600_ _1220_ _1237_ _1549_ VPWR VGND sg13g2_nor2_2
X_5580_ net255 VGND VPWR net488 falu_i.falutop.div_inst.a\[3\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_2792_ _2146_ net542 VPWR VGND sg13g2_inv_2
XFILLER_7_360 VPWR VGND sg13g2_fill_1
X_4531_ _1479_ _1480_ _1309_ _1481_ VPWR VGND sg13g2_nand3_1
XFILLER_11_1007 VPWR VGND sg13g2_decap_8
X_4462_ net765 net736 net566 _1413_ VPWR VGND sg13g2_mux2_1
Xhold316 _0332_ VPWR VGND net968 sg13g2_dlygate4sd3_1
Xhold305 ppwm_i.u_ppwm.u_mem.memory\[91\] VPWR VGND net957 sg13g2_dlygate4sd3_1
Xhold338 _0454_ VPWR VGND net990 sg13g2_dlygate4sd3_1
Xhold327 _0266_ VPWR VGND net979 sg13g2_dlygate4sd3_1
Xhold349 falu_i.falutop.i2c_inst.state\[1\] VPWR VGND net1001 sg13g2_dlygate4sd3_1
X_3413_ _2251_ ppwm_i.u_ppwm.global_counter\[10\] _0590_ _0591_ VPWR VGND sg13g2_nor3_1
X_4393_ VPWR VGND _1301_ _1345_ _1299_ net616 _1346_ _1283_ sg13g2_a221oi_1
Xfanout807 net808 net807 VPWR VGND sg13g2_buf_8
Xfanout829 net830 net829 VPWR VGND sg13g2_buf_8
Xfanout818 net820 net818 VPWR VGND sg13g2_buf_8
X_3344_ VPWR VGND _0520_ _0521_ _0519_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] _0522_
+ _2250_ sg13g2_a221oi_1
X_3275_ net812 VPWR _0459_ VGND _2258_ _0457_ sg13g2_o21ai_1
X_5014_ _1955_ _1946_ _1956_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_275 VPWR VGND sg13g2_decap_8
XFILLER_27_938 VPWR VGND sg13g2_decap_8
XFILLER_34_481 VPWR VGND sg13g2_fill_1
XFILLER_10_838 VPWR VGND sg13g2_decap_8
XFILLER_21_164 VPWR VGND sg13g2_fill_1
X_4729_ _1675_ VPWR _1676_ VGND _1374_ _1670_ sg13g2_o21ai_1
XFILLER_1_514 VPWR VGND sg13g2_decap_8
XFILLER_18_949 VPWR VGND sg13g2_decap_8
XFILLER_44_278 VPWR VGND sg13g2_decap_4
XFILLER_26_993 VPWR VGND sg13g2_decap_8
XFILLER_41_941 VPWR VGND sg13g2_decap_8
XFILLER_16_83 VPWR VGND sg13g2_decap_8
XFILLER_25_492 VPWR VGND sg13g2_fill_1
XFILLER_13_665 VPWR VGND sg13g2_decap_4
XFILLER_34_1018 VPWR VGND sg13g2_decap_8
XFILLER_40_495 VPWR VGND sg13g2_fill_1
XFILLER_5_820 VPWR VGND sg13g2_fill_1
XFILLER_5_853 VPWR VGND sg13g2_decap_8
XFILLER_4_363 VPWR VGND sg13g2_fill_2
X_3060_ _2412_ _2413_ _2411_ _2414_ VPWR VGND sg13g2_nand3_1
XFILLER_17_960 VPWR VGND sg13g2_decap_8
XFILLER_35_278 VPWR VGND sg13g2_decap_8
X_3962_ VGND VPWR _2164_ net672 _0200_ _1009_ sg13g2_a21oi_1
X_3893_ net839 VPWR _0975_ VGND ppwm_i.u_ppwm.u_mem.memory\[66\] net676 sg13g2_o21ai_1
X_2913_ _2267_ net553 VPWR VGND sg13g2_inv_2
X_2844_ VPWR _2198_ net443 VGND sg13g2_inv_1
XFILLER_32_996 VPWR VGND sg13g2_decap_8
X_5563_ net124 VGND VPWR _0322_ falu_i.falutop.alu_data_in\[9\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_2
X_4514_ _1464_ net743 net710 VPWR VGND sg13g2_nand2_1
Xhold102 ppwm_i.u_ppwm.u_mem.memory\[62\] VPWR VGND net474 sg13g2_dlygate4sd3_1
Xhold113 falu_i.falutop.div_inst.acc\[7\] VPWR VGND net485 sg13g2_dlygate4sd3_1
X_5494_ net291 VGND VPWR net919 falu_i.falutop.div_inst.i\[1\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
Xhold124 ppwm_i.u_ppwm.u_mem.memory\[15\] VPWR VGND net496 sg13g2_dlygate4sd3_1
Xhold135 _0025_ VPWR VGND net507 sg13g2_dlygate4sd3_1
X_4445_ _1395_ _1396_ _1397_ VPWR VGND sg13g2_nor2_1
Xhold168 ppwm_i.u_ppwm.u_mem.memory\[108\] VPWR VGND net540 sg13g2_dlygate4sd3_1
Xhold157 _0205_ VPWR VGND net529 sg13g2_dlygate4sd3_1
Xhold146 ppwm_i.u_ppwm.u_mem.memory\[87\] VPWR VGND net518 sg13g2_dlygate4sd3_1
Xhold179 ppwm_i.u_ppwm.u_mem.memory\[78\] VPWR VGND net551 sg13g2_dlygate4sd3_1
Xfanout604 _2374_ net604 VPWR VGND sg13g2_buf_8
Xfanout615 _1317_ net615 VPWR VGND sg13g2_buf_8
X_4376_ _1259_ _1302_ _1329_ VPWR VGND sg13g2_nor2b_1
X_3327_ _0506_ _2308_ _0505_ VPWR VGND sg13g2_nand2_1
Xfanout637 _1134_ net637 VPWR VGND sg13g2_buf_8
Xfanout626 _1077_ net626 VPWR VGND sg13g2_buf_8
Xfanout648 net650 net648 VPWR VGND sg13g2_buf_8
Xfanout659 net663 net659 VPWR VGND sg13g2_buf_8
XFILLER_39_551 VPWR VGND sg13g2_fill_1
X_3258_ net796 net1130 _0058_ VPWR VGND sg13g2_nor2_1
XFILLER_2_1027 VPWR VGND sg13g2_fill_2
XFILLER_2_1016 VPWR VGND sg13g2_decap_8
X_3189_ net1117 _0400_ _0402_ VPWR VGND sg13g2_and2_1
XFILLER_42_727 VPWR VGND sg13g2_fill_2
XFILLER_26_278 VPWR VGND sg13g2_fill_2
XFILLER_23_996 VPWR VGND sg13g2_decap_8
XFILLER_2_834 VPWR VGND sg13g2_decap_8
XFILLER_2_801 VPWR VGND sg13g2_fill_2
XFILLER_49_304 VPWR VGND sg13g2_fill_1
XFILLER_49_326 VPWR VGND sg13g2_decap_8
XFILLER_18_702 VPWR VGND sg13g2_fill_1
XFILLER_45_510 VPWR VGND sg13g2_decap_4
XFILLER_18_713 VPWR VGND sg13g2_decap_8
XFILLER_45_543 VPWR VGND sg13g2_decap_8
XFILLER_9_400 VPWR VGND sg13g2_decap_4
XFILLER_14_985 VPWR VGND sg13g2_decap_8
X_4230_ VGND VPWR net781 falu_i.falutop.div_inst.a\[3\] _1195_ _1194_ sg13g2_a21oi_1
X_4161_ net568 net633 _1145_ VPWR VGND sg13g2_nor2b_1
X_4092_ falu_i.falutop.div_inst.i\[1\] net525 net409 _1095_ VPWR VGND sg13g2_nand3_1
X_3112_ net817 VPWR _0352_ VGND net881 net988 sg13g2_o21ai_1
X_3043_ VGND VPWR _2395_ _2396_ _2397_ _2254_ sg13g2_a21oi_1
X_4994_ _1903_ VPWR _1936_ VGND _1215_ _1904_ sg13g2_o21ai_1
XFILLER_23_215 VPWR VGND sg13g2_decap_4
XFILLER_17_1002 VPWR VGND sg13g2_decap_8
X_3945_ net837 VPWR _1001_ VGND net401 net648 sg13g2_o21ai_1
XFILLER_20_944 VPWR VGND sg13g2_decap_8
XFILLER_23_29 VPWR VGND sg13g2_decap_8
X_3876_ VGND VPWR _2195_ net671 _0157_ _0966_ sg13g2_a21oi_1
X_2827_ VPWR _2181_ net843 VGND sg13g2_inv_1
X_5546_ net313 VGND VPWR net1063 falu_i.falutop.i2c_inst.result\[10\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_5477_ net331 VGND VPWR net874 falu_i.falutop.data_in\[8\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_4428_ _1380_ net766 net745 net769 net741 VPWR VGND sg13g2_a22oi_1
X_4359_ _1309_ _1311_ _1308_ _1312_ VPWR VGND sg13g2_nand3_1
XFILLER_47_819 VPWR VGND sg13g2_fill_1
XFILLER_24_1028 VPWR VGND sg13g2_fill_1
XFILLER_27_554 VPWR VGND sg13g2_fill_1
XFILLER_42_524 VPWR VGND sg13g2_fill_2
XFILLER_27_598 VPWR VGND sg13g2_decap_4
XFILLER_23_793 VPWR VGND sg13g2_decap_8
XFILLER_10_443 VPWR VGND sg13g2_decap_8
XFILLER_11_944 VPWR VGND sg13g2_decap_8
XFILLER_13_40 VPWR VGND sg13g2_fill_2
XFILLER_7_937 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_1
XFILLER_46_841 VPWR VGND sg13g2_fill_1
XFILLER_45_351 VPWR VGND sg13g2_decap_8
X_3730_ net575 VPWR _0888_ VGND _0884_ _0886_ sg13g2_o21ai_1
X_3661_ _0824_ _0825_ _0826_ VPWR VGND sg13g2_and2_1
X_3592_ net577 VPWR _0762_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] net588 sg13g2_o21ai_1
X_5400_ net252 VGND VPWR _0159_ ppwm_i.u_ppwm.u_mem.memory\[59\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_5331_ net39 VGND VPWR net1195 ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_1
X_5262_ net172 VGND VPWR net382 ppwm_i.u_ppwm.u_pwm.cmp_value\[0\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
X_4213_ _1182_ net567 _1181_ _1131_ _2290_ VPWR VGND sg13g2_a22oi_1
X_5193_ _2111_ net777 falu_i.falutop.data_in\[0\] VPWR VGND sg13g2_nand2_1
X_4144_ _0252_ net526 _1096_ _1138_ _1095_ VPWR VGND sg13g2_a22oi_1
XFILLER_49_690 VPWR VGND sg13g2_decap_8
X_4075_ falu_i.falutop.i2c_inst.result\[10\] _0343_ _1079_ VPWR VGND sg13g2_and2_1
X_3026_ VPWR VGND _2187_ net789 net690 _2192_ _2380_ net697 sg13g2_a221oi_1
XFILLER_37_863 VPWR VGND sg13g2_decap_8
X_4977_ _1918_ _1890_ _1920_ VPWR VGND sg13g2_xor2_1
X_5352__348 VPWR VGND net348 sg13g2_tiehi
Xclkload5 clknet_leaf_35_clk clkload5/Y VPWR VGND sg13g2_inv_4
X_3928_ VGND VPWR _2175_ net674 _0183_ _0992_ sg13g2_a21oi_1
X_3859_ net829 VPWR _0958_ VGND net434 net664 sg13g2_o21ai_1
XFILLER_30_1021 VPWR VGND sg13g2_decap_8
XFILLER_4_929 VPWR VGND sg13g2_decap_8
X_5529_ net153 VGND VPWR net490 falu_i.falutop.div_inst.acc\[2\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_8_1000 VPWR VGND sg13g2_decap_8
XFILLER_15_502 VPWR VGND sg13g2_fill_2
XFILLER_28_863 VPWR VGND sg13g2_decap_4
XFILLER_15_579 VPWR VGND sg13g2_decap_8
XFILLER_11_752 VPWR VGND sg13g2_fill_2
XFILLER_24_61 VPWR VGND sg13g2_fill_2
XFILLER_7_756 VPWR VGND sg13g2_fill_1
XFILLER_3_973 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_46_660 VPWR VGND sg13g2_fill_1
XFILLER_19_863 VPWR VGND sg13g2_decap_8
X_4900_ _1805_ VPWR _1844_ VGND _1801_ _1802_ sg13g2_o21ai_1
X_4831_ _1777_ _1776_ _1708_ VPWR VGND sg13g2_nand2b_1
X_5258__179 VPWR VGND net179 sg13g2_tiehi
X_4762_ _1707_ _1681_ _1709_ VPWR VGND sg13g2_xor2_1
X_3713_ _0759_ net569 _0872_ _0873_ VPWR VGND sg13g2_nor3_1
XFILLER_14_1027 VPWR VGND sg13g2_fill_2
X_4693_ _1640_ _1567_ _1641_ VPWR VGND sg13g2_xor2_1
X_3644_ _0809_ _0810_ _0081_ VPWR VGND sg13g2_nor2_1
X_3575_ VPWR VGND _0745_ net799 _0732_ _2247_ _0077_ net572 sg13g2_a221oi_1
X_5314_ net73 VGND VPWR net1197 ppwm_i.u_ppwm.pwm_value\[1\] clknet_leaf_19_clk sg13g2_dfrbpq_1
X_5245_ net205 VGND VPWR _0007_ falu_i.falutop.i2c_inst.data_in\[3\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
Xhold28 _0280_ VPWR VGND net400 sg13g2_dlygate4sd3_1
Xhold17 _0337_ VPWR VGND net389 sg13g2_dlygate4sd3_1
X_5176_ VGND VPWR _2305_ net619 _0318_ _2105_ sg13g2_a21oi_1
Xhold39 falu_i.falutop.div_inst.quo\[2\] VPWR VGND net411 sg13g2_dlygate4sd3_1
X_4127_ VGND VPWR _1127_ _1128_ _1129_ _1111_ sg13g2_a21oi_1
X_4058_ net380 net622 _0227_ VPWR VGND sg13g2_nor2_1
X_3009_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[97\] net709 net690 ppwm_i.u_ppwm.u_mem.memory\[104\]
+ _2363_ net694 sg13g2_a221oi_1
XFILLER_25_855 VPWR VGND sg13g2_decap_8
XFILLER_40_825 VPWR VGND sg13g2_fill_2
XFILLER_40_858 VPWR VGND sg13g2_decap_4
XFILLER_3_269 VPWR VGND sg13g2_fill_2
XFILLER_3_247 VPWR VGND sg13g2_decap_4
XFILLER_0_932 VPWR VGND sg13g2_decap_8
XFILLER_48_914 VPWR VGND sg13g2_decap_8
XFILLER_19_115 VPWR VGND sg13g2_fill_1
XFILLER_16_811 VPWR VGND sg13g2_fill_1
XFILLER_15_332 VPWR VGND sg13g2_decap_8
XFILLER_37_1027 VPWR VGND sg13g2_fill_2
XFILLER_16_888 VPWR VGND sg13g2_decap_8
XFILLER_7_542 VPWR VGND sg13g2_fill_1
Xhold509 _0091_ VPWR VGND net1161 sg13g2_dlygate4sd3_1
XFILLER_7_553 VPWR VGND sg13g2_decap_4
X_3360_ VPWR VGND ppwm_i.u_ppwm.pwm_value\[2\] _0537_ _2272_ ppwm_i.u_ppwm.pwm_value\[3\]
+ _0538_ _2271_ sg13g2_a221oi_1
X_3291_ VGND VPWR _2273_ ppwm_i.u_ppwm.u_pwm.cmp_value\[9\] _0474_ _0473_ sg13g2_a21oi_1
X_5030_ _1590_ VPWR _1972_ VGND _1968_ _1971_ sg13g2_o21ai_1
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_22_803 VPWR VGND sg13g2_decap_8
X_4814_ _1760_ net728 falu_i.falutop.alu_data_in\[7\] net755 VPWR VGND sg13g2_and3_1
X_5271__154 VPWR VGND net154 sg13g2_tiehi
X_4745_ _1629_ VPWR _1692_ VGND _1392_ _1630_ sg13g2_o21ai_1
XFILLER_21_379 VPWR VGND sg13g2_decap_4
X_4676_ _1624_ net753 net741 net768 net723 VPWR VGND sg13g2_a22oi_1
X_3627_ net580 VPWR _0795_ VGND net783 net589 sg13g2_o21ai_1
X_3558_ _0729_ _2247_ net600 VPWR VGND sg13g2_xnor2_1
XFILLER_0_206 VPWR VGND sg13g2_fill_1
X_3489_ VGND VPWR net589 _0662_ _0664_ _0663_ sg13g2_a21oi_1
XFILLER_5_1014 VPWR VGND sg13g2_decap_8
X_5228_ VGND VPWR net625 _2136_ _0339_ _2135_ sg13g2_a21oi_1
X_5159_ VPWR _0311_ net953 VGND sg13g2_inv_1
XFILLER_29_468 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_decap_4
Xclkbuf_leaf_36_clk clknet_3_5__leaf_clk clknet_leaf_36_clk VPWR VGND sg13g2_buf_8
XFILLER_40_600 VPWR VGND sg13g2_decap_8
XFILLER_40_622 VPWR VGND sg13g2_decap_8
XFILLER_9_807 VPWR VGND sg13g2_decap_4
XFILLER_4_534 VPWR VGND sg13g2_fill_1
XFILLER_47_232 VPWR VGND sg13g2_fill_1
XFILLER_29_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_27_clk clknet_3_6__leaf_clk clknet_leaf_27_clk VPWR VGND sg13g2_buf_8
XFILLER_16_630 VPWR VGND sg13g2_fill_2
XFILLER_44_972 VPWR VGND sg13g2_decap_8
XFILLER_15_140 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_fill_2
X_2860_ VPWR _2214_ net845 VGND sg13g2_inv_1
XFILLER_7_350 VPWR VGND sg13g2_fill_2
X_4530_ _1480_ _1477_ _1478_ VPWR VGND sg13g2_nand2_1
Xhold317 ppwm_i.u_ppwm.u_mem.memory\[42\] VPWR VGND net969 sg13g2_dlygate4sd3_1
XFILLER_8_895 VPWR VGND sg13g2_decap_8
X_4461_ _1409_ _1411_ _1261_ _1412_ VPWR VGND sg13g2_nand3_1
Xhold306 _0190_ VPWR VGND net958 sg13g2_dlygate4sd3_1
Xhold339 _0062_ VPWR VGND net991 sg13g2_dlygate4sd3_1
X_3412_ net784 _2266_ _0590_ VPWR VGND sg13g2_nor2_1
Xhold328 ppwm_i.u_ppwm.u_ex.state_q\[0\] VPWR VGND net980 sg13g2_dlygate4sd3_1
X_4392_ _1320_ _1328_ _1316_ _1345_ VPWR VGND _1344_ sg13g2_nand4_1
Xfanout819 net820 net819 VPWR VGND sg13g2_buf_2
Xfanout808 net811 net808 VPWR VGND sg13g2_buf_8
X_3343_ _2242_ net784 _0521_ VPWR VGND sg13g2_nor2_1
X_3274_ VGND VPWR _2259_ _0455_ _0063_ _0458_ sg13g2_a21oi_1
X_5013_ _1955_ _1948_ _1953_ VPWR VGND sg13g2_xnor2_1
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_38_298 VPWR VGND sg13g2_fill_1
XFILLER_26_438 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_18_clk clknet_3_4__leaf_clk clknet_leaf_18_clk VPWR VGND sg13g2_buf_8
XFILLER_19_490 VPWR VGND sg13g2_fill_2
XFILLER_41_408 VPWR VGND sg13g2_decap_4
XFILLER_34_493 VPWR VGND sg13g2_decap_8
X_2989_ VPWR VGND _2342_ net787 _2341_ _2339_ _2343_ _2340_ sg13g2_a221oi_1
X_4728_ VPWR VGND _1247_ _1674_ _1671_ _1244_ _1675_ _1327_ sg13g2_a221oi_1
X_4659_ net750 net565 _1607_ VPWR VGND sg13g2_nor2_1
XFILLER_27_1015 VPWR VGND sg13g2_decap_8
X_5505__265 VPWR VGND net265 sg13g2_tiehi
XFILLER_18_928 VPWR VGND sg13g2_decap_8
XFILLER_17_449 VPWR VGND sg13g2_decap_8
XFILLER_26_972 VPWR VGND sg13g2_decap_8
XFILLER_32_408 VPWR VGND sg13g2_decap_4
XFILLER_13_633 VPWR VGND sg13g2_fill_1
XFILLER_16_73 VPWR VGND sg13g2_decap_4
XFILLER_12_154 VPWR VGND sg13g2_decap_4
XFILLER_41_997 VPWR VGND sg13g2_decap_8
XFILLER_9_648 VPWR VGND sg13g2_decap_8
XFILLER_5_832 VPWR VGND sg13g2_decap_8
XFILLER_4_386 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_0_592 VPWR VGND sg13g2_fill_2
XFILLER_36_725 VPWR VGND sg13g2_decap_8
XFILLER_16_460 VPWR VGND sg13g2_decap_4
X_3961_ net838 VPWR _1009_ VGND ppwm_i.u_ppwm.u_mem.memory\[100\] net672 sg13g2_o21ai_1
X_2912_ _2266_ ppwm_i.u_ppwm.global_counter\[11\] VPWR VGND sg13g2_inv_2
X_3892_ VGND VPWR _2189_ net669 _0165_ _0974_ sg13g2_a21oi_1
XFILLER_32_975 VPWR VGND sg13g2_decap_8
X_2843_ VPWR _2197_ net469 VGND sg13g2_inv_1
X_5562_ net133 VGND VPWR net1159 falu_i.falutop.alu_data_in\[8\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_4513_ _1421_ VPWR _1463_ VGND _1393_ _1419_ sg13g2_o21ai_1
Xhold103 falu_i.falutop.div_inst.a\[2\] VPWR VGND net475 sg13g2_dlygate4sd3_1
Xhold114 _0293_ VPWR VGND net486 sg13g2_dlygate4sd3_1
X_5493_ net295 VGND VPWR net527 falu_i.falutop.div_inst.i\[0\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
Xhold125 _0114_ VPWR VGND net497 sg13g2_dlygate4sd3_1
Xhold158 ppwm_i.u_ppwm.u_mem.memory\[46\] VPWR VGND net530 sg13g2_dlygate4sd3_1
X_4444_ _1396_ net744 net721 VPWR VGND sg13g2_nand2_1
Xclkbuf_leaf_7_clk clknet_3_5__leaf_clk clknet_leaf_7_clk VPWR VGND sg13g2_buf_8
Xhold136 ppwm_i.u_ppwm.u_mem.memory\[26\] VPWR VGND net508 sg13g2_dlygate4sd3_1
Xhold147 _0187_ VPWR VGND net519 sg13g2_dlygate4sd3_1
Xfanout605 net606 net605 VPWR VGND sg13g2_buf_8
X_4375_ VPWR VGND _1220_ net640 _1327_ _1223_ _1328_ _1326_ sg13g2_a221oi_1
Xhold169 ppwm_i.u_ppwm.u_mem.memory\[88\] VPWR VGND net541 sg13g2_dlygate4sd3_1
Xfanout649 net650 net649 VPWR VGND sg13g2_buf_8
X_3326_ _2254_ VPWR _0505_ VGND net708 _2307_ sg13g2_o21ai_1
Xfanout638 net640 net638 VPWR VGND sg13g2_buf_8
Xfanout627 net629 net627 VPWR VGND sg13g2_buf_8
Xfanout616 _1281_ net616 VPWR VGND sg13g2_buf_8
X_3257_ _0447_ net1129 _0445_ VPWR VGND sg13g2_xnor2_1
X_3188_ _0400_ net1112 _0034_ VPWR VGND sg13g2_nor2_1
XFILLER_22_452 VPWR VGND sg13g2_fill_2
XFILLER_23_975 VPWR VGND sg13g2_decap_8
XFILLER_10_625 VPWR VGND sg13g2_decap_8
XFILLER_2_813 VPWR VGND sg13g2_decap_8
X_5362__328 VPWR VGND net328 sg13g2_tiehi
XFILLER_40_1023 VPWR VGND sg13g2_decap_4
XFILLER_45_533 VPWR VGND sg13g2_fill_2
XFILLER_17_224 VPWR VGND sg13g2_decap_8
XFILLER_18_769 VPWR VGND sg13g2_fill_2
XFILLER_13_441 VPWR VGND sg13g2_decap_8
XFILLER_13_452 VPWR VGND sg13g2_fill_1
XFILLER_14_964 VPWR VGND sg13g2_decap_8
XFILLER_25_290 VPWR VGND sg13g2_fill_2
XFILLER_43_71 VPWR VGND sg13g2_decap_4
XFILLER_9_434 VPWR VGND sg13g2_decap_8
XFILLER_9_467 VPWR VGND sg13g2_fill_2
XFILLER_5_684 VPWR VGND sg13g2_decap_8
X_5408__236 VPWR VGND net236 sg13g2_tiehi
X_4160_ net797 net607 _0263_ VPWR VGND sg13g2_nor2_1
X_3111_ _2439_ net987 _0351_ VPWR VGND sg13g2_nor2_1
X_4091_ _1093_ net997 _0244_ VPWR VGND sg13g2_nor2_1
XFILLER_49_894 VPWR VGND sg13g2_decap_8
X_3042_ VPWR VGND _2194_ net790 net697 _2178_ _2396_ net703 sg13g2_a221oi_1
X_4993_ _1913_ VPWR _1935_ VGND _1901_ _1914_ sg13g2_o21ai_1
XFILLER_24_739 VPWR VGND sg13g2_decap_8
X_3944_ VGND VPWR _2170_ net673 _0191_ _1000_ sg13g2_a21oi_1
X_3875_ net835 VPWR _0966_ VGND ppwm_i.u_ppwm.u_mem.memory\[57\] net671 sg13g2_o21ai_1
XFILLER_20_923 VPWR VGND sg13g2_decap_8
X_2826_ VPWR _2180_ net551 VGND sg13g2_inv_1
X_5545_ net355 VGND VPWR net1065 falu_i.falutop.i2c_inst.result\[9\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_5476_ net333 VGND VPWR net872 falu_i.falutop.data_in\[7\] clknet_leaf_2_clk sg13g2_dfrbpq_2
X_4427_ VPWR _1379_ _1378_ VGND sg13g2_inv_1
X_5316__69 VPWR VGND net69 sg13g2_tiehi
X_5331__39 VPWR VGND net39 sg13g2_tiehi
X_4358_ VGND VPWR _1311_ net770 net726 sg13g2_or2_1
XFILLER_47_809 VPWR VGND sg13g2_fill_2
X_3309_ _0490_ _0489_ _2422_ VPWR VGND sg13g2_nand2b_1
X_4289_ _1242_ _1241_ VPWR VGND _1240_ sg13g2_nand2b_2
XFILLER_15_706 VPWR VGND sg13g2_fill_1
XFILLER_27_577 VPWR VGND sg13g2_decap_8
XFILLER_10_400 VPWR VGND sg13g2_fill_1
XFILLER_11_923 VPWR VGND sg13g2_decap_8
XFILLER_23_772 VPWR VGND sg13g2_decap_8
XFILLER_7_916 VPWR VGND sg13g2_decap_8
XFILLER_6_415 VPWR VGND sg13g2_decap_4
XFILLER_10_477 VPWR VGND sg13g2_decap_4
XFILLER_18_599 VPWR VGND sg13g2_fill_1
XFILLER_14_761 VPWR VGND sg13g2_fill_1
X_3660_ VGND VPWR _0815_ _0823_ _0825_ _0618_ sg13g2_a21oi_1
X_3591_ VGND VPWR ppwm_i.u_ppwm.global_counter\[16\] net592 _0761_ _0760_ sg13g2_a21oi_1
XFILLER_9_297 VPWR VGND sg13g2_decap_4
X_5330_ net41 VGND VPWR net1170 ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_2
XFILLER_5_470 VPWR VGND sg13g2_decap_8
X_5261_ net173 VGND VPWR _0023_ ppwm_i.u_ppwm.u_mem.data_sync2 clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
X_4212_ _1181_ _1110_ _1129_ VPWR VGND sg13g2_xnor2_1
X_5192_ _2110_ net413 net622 VPWR VGND sg13g2_nand2_1
X_4143_ _1139_ net525 net778 VPWR VGND sg13g2_nand2b_1
X_4074_ net908 net775 net684 _0243_ VPWR VGND sg13g2_mux2_1
X_3025_ _2379_ net694 _2182_ net703 _2176_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_831 VPWR VGND sg13g2_decap_8
XFILLER_36_363 VPWR VGND sg13g2_fill_2
X_4976_ _1918_ _1890_ _1919_ VPWR VGND sg13g2_nor2b_1
X_3927_ net841 VPWR _0992_ VGND net930 net674 sg13g2_o21ai_1
X_3858_ VGND VPWR _2201_ net658 _0148_ _0957_ sg13g2_a21oi_1
Xclkload6 clkload6/Y clknet_leaf_36_clk VPWR VGND sg13g2_inv_8
XFILLER_30_1000 VPWR VGND sg13g2_decap_8
XFILLER_4_908 VPWR VGND sg13g2_decap_8
X_2809_ VPWR _2163_ net539 VGND sg13g2_inv_1
X_3789_ net828 VPWR _0923_ VGND ppwm_i.u_ppwm.u_mem.memory\[14\] net661 sg13g2_o21ai_1
X_5528_ net161 VGND VPWR net499 falu_i.falutop.div_inst.acc\[1\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_5459_ net50 VGND VPWR net514 ppwm_i.u_ppwm.u_mem.bit_count\[6\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_1
X_5281__134 VPWR VGND net134 sg13g2_tiehi
X_5426__188 VPWR VGND net188 sg13g2_tiehi
X_5458__54 VPWR VGND net54 sg13g2_tiehi
XFILLER_28_820 VPWR VGND sg13g2_fill_2
XFILLER_42_333 VPWR VGND sg13g2_decap_8
XFILLER_23_580 VPWR VGND sg13g2_fill_1
X_5433__159 VPWR VGND net159 sg13g2_tiehi
XFILLER_7_713 VPWR VGND sg13g2_decap_4
XFILLER_6_201 VPWR VGND sg13g2_decap_4
XFILLER_10_274 VPWR VGND sg13g2_fill_1
XFILLER_3_952 VPWR VGND sg13g2_decap_8
XFILLER_2_484 VPWR VGND sg13g2_decap_8
XFILLER_34_8 VPWR VGND sg13g2_fill_1
XFILLER_49_81 VPWR VGND sg13g2_fill_1
X_5303__94 VPWR VGND net94 sg13g2_tiehi
XFILLER_37_105 VPWR VGND sg13g2_decap_4
X_5520__198 VPWR VGND net198 sg13g2_tiehi
XFILLER_19_842 VPWR VGND sg13g2_decap_8
XFILLER_1_99 VPWR VGND sg13g2_decap_4
XFILLER_18_374 VPWR VGND sg13g2_decap_8
X_4830_ _1775_ _1684_ _1776_ VPWR VGND sg13g2_xor2_1
XFILLER_14_591 VPWR VGND sg13g2_fill_2
X_4761_ _1708_ _1681_ _1707_ VPWR VGND sg13g2_nand2b_1
X_3712_ VGND VPWR net581 _0761_ _0872_ _0871_ sg13g2_a21oi_1
XFILLER_14_1006 VPWR VGND sg13g2_decap_8
X_4692_ _1640_ _1638_ _1639_ VPWR VGND sg13g2_xnor2_1
X_3643_ net821 VPWR _0810_ VGND net1167 _0614_ sg13g2_o21ai_1
X_3574_ _0740_ _0744_ _0745_ VPWR VGND sg13g2_and2_1
X_5313_ net75 VGND VPWR _0072_ ppwm_i.u_ppwm.pwm_value\[0\] clknet_leaf_19_clk sg13g2_dfrbpq_2
X_5244_ net207 VGND VPWR _0006_ falu_i.falutop.i2c_inst.data_in\[2\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_5175_ net1153 net619 _2105_ VPWR VGND sg13g2_nor2_1
Xhold18 ppwm_i.u_ppwm.u_mem.memory\[92\] VPWR VGND net390 sg13g2_dlygate4sd3_1
Xhold29 ppwm_i.u_ppwm.u_mem.memory\[93\] VPWR VGND net401 sg13g2_dlygate4sd3_1
X_4126_ _1128_ falu_i.falutop.div_inst.b1\[6\] falu_i.falutop.div_inst.acc\[6\] VPWR
+ VGND sg13g2_xnor2_1
XFILLER_44_609 VPWR VGND sg13g2_decap_4
X_4057_ _1078_ net815 net638 VPWR VGND sg13g2_nand2_2
X_3008_ _2362_ net697 ppwm_i.u_ppwm.u_mem.memory\[90\] net702 ppwm_i.u_ppwm.u_mem.memory\[111\]
+ VPWR VGND sg13g2_a22oi_1
X_4959_ _1863_ VPWR _1902_ VGND _1856_ _1864_ sg13g2_o21ai_1
XFILLER_0_911 VPWR VGND sg13g2_decap_8
XFILLER_0_988 VPWR VGND sg13g2_decap_8
X_5300__97 VPWR VGND net97 sg13g2_tiehi
XFILLER_43_620 VPWR VGND sg13g2_fill_1
XFILLER_43_631 VPWR VGND sg13g2_decap_4
XFILLER_37_1006 VPWR VGND sg13g2_decap_8
XFILLER_16_867 VPWR VGND sg13g2_decap_8
XFILLER_27_193 VPWR VGND sg13g2_decap_8
XFILLER_30_358 VPWR VGND sg13g2_fill_1
X_3290_ VPWR VGND ppwm_i.u_ppwm.u_pwm.counter\[8\] _0472_ _2280_ ppwm_i.u_ppwm.u_pwm.counter\[9\]
+ _0473_ _2279_ sg13g2_a221oi_1
XFILLER_3_771 VPWR VGND sg13g2_fill_1
XFILLER_3_760 VPWR VGND sg13g2_fill_1
XFILLER_25_4 VPWR VGND sg13g2_fill_1
XFILLER_39_959 VPWR VGND sg13g2_decap_8
XFILLER_19_650 VPWR VGND sg13g2_decap_8
XFILLER_20_1021 VPWR VGND sg13g2_decap_8
XFILLER_26_609 VPWR VGND sg13g2_decap_4
XFILLER_47_981 VPWR VGND sg13g2_decap_8
XFILLER_25_119 VPWR VGND sg13g2_fill_2
XFILLER_33_152 VPWR VGND sg13g2_fill_1
X_4813_ _1759_ net723 net761 VPWR VGND sg13g2_nand2_1
XFILLER_22_859 VPWR VGND sg13g2_decap_8
X_4744_ _1690_ _1687_ _1691_ VPWR VGND sg13g2_xor2_1
XFILLER_30_870 VPWR VGND sg13g2_fill_1
X_4675_ _2295_ _2301_ _1622_ _1623_ VPWR VGND sg13g2_nor3_1
X_3626_ VPWR _0794_ _0793_ VGND sg13g2_inv_1
X_3557_ _0727_ _0728_ _0076_ VPWR VGND sg13g2_nor2_1
XFILLER_0_218 VPWR VGND sg13g2_decap_8
X_5227_ _2136_ falu_i.falutop.data_in\[11\] _2134_ VPWR VGND sg13g2_xnor2_1
X_3488_ net579 VPWR _0663_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] net589 sg13g2_o21ai_1
X_5158_ _2095_ _2094_ net774 _1078_ net952 VPWR VGND sg13g2_a22oi_1
XFILLER_29_425 VPWR VGND sg13g2_fill_1
XFILLER_45_929 VPWR VGND sg13g2_decap_8
X_4109_ falu_i.falutop.div_inst.b1\[6\] falu_i.falutop.div_inst.acc\[6\] _1111_ VPWR
+ VGND sg13g2_nor2b_1
X_5089_ _2026_ _2028_ _2029_ VPWR VGND sg13g2_nor2_1
XFILLER_38_981 VPWR VGND sg13g2_decap_8
XFILLER_13_815 VPWR VGND sg13g2_fill_1
XFILLER_13_859 VPWR VGND sg13g2_decap_8
XFILLER_24_185 VPWR VGND sg13g2_fill_1
X_5451__82 VPWR VGND net82 sg13g2_tiehi
XFILLER_4_513 VPWR VGND sg13g2_fill_2
XFILLER_43_1010 VPWR VGND sg13g2_decap_8
XFILLER_48_723 VPWR VGND sg13g2_fill_1
XFILLER_47_211 VPWR VGND sg13g2_fill_1
XFILLER_0_785 VPWR VGND sg13g2_decap_8
X_5341__370 VPWR VGND net370 sg13g2_tiehi
XFILLER_47_266 VPWR VGND sg13g2_fill_2
XFILLER_29_970 VPWR VGND sg13g2_decap_8
XFILLER_44_951 VPWR VGND sg13g2_decap_8
XFILLER_35_439 VPWR VGND sg13g2_decap_4
X_5372__308 VPWR VGND net308 sg13g2_tiehi
XFILLER_43_450 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_fill_1
XFILLER_30_133 VPWR VGND sg13g2_fill_2
XFILLER_12_881 VPWR VGND sg13g2_decap_8
XFILLER_8_874 VPWR VGND sg13g2_decap_8
Xhold307 ppwm_i.u_ppwm.u_mem.memory\[28\] VPWR VGND net959 sg13g2_dlygate4sd3_1
X_4460_ _1356_ _1358_ _1353_ _1411_ VPWR VGND sg13g2_nand3_1
X_3411_ VGND VPWR _2243_ ppwm_i.u_ppwm.global_counter\[19\] _0589_ net591 sg13g2_a21oi_1
Xhold318 _0141_ VPWR VGND net970 sg13g2_dlygate4sd3_1
X_4391_ _1344_ _1338_ _1343_ _1336_ _1329_ VPWR VGND sg13g2_a22oi_1
Xhold329 _2425_ VPWR VGND net981 sg13g2_dlygate4sd3_1
X_3342_ ppwm_i.u_ppwm.pwm_value\[0\] ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] _0520_ VPWR
+ VGND sg13g2_nor2b_1
Xfanout809 net811 net809 VPWR VGND sg13g2_buf_8
X_3273_ _0458_ net813 _0457_ VPWR VGND sg13g2_nand2_1
XFILLER_39_701 VPWR VGND sg13g2_decap_8
XFILLER_39_712 VPWR VGND sg13g2_fill_1
X_5012_ _1948_ _1953_ _1954_ VPWR VGND sg13g2_nor2_1
XFILLER_38_255 VPWR VGND sg13g2_fill_1
X_5418__216 VPWR VGND net216 sg13g2_tiehi
X_5533__120 VPWR VGND net120 sg13g2_tiehi
XFILLER_35_984 VPWR VGND sg13g2_decap_8
XFILLER_22_656 VPWR VGND sg13g2_fill_1
X_2988_ VPWR VGND _2210_ net708 net688 _2201_ _2342_ net701 sg13g2_a221oi_1
XFILLER_21_155 VPWR VGND sg13g2_fill_1
X_4727_ _1673_ VPWR _1674_ VGND _1245_ _1672_ sg13g2_o21ai_1
X_4658_ _1606_ _1309_ _1605_ VPWR VGND sg13g2_nand2_1
X_3609_ VGND VPWR net590 _0776_ _0778_ _0777_ sg13g2_a21oi_1
X_4589_ _1472_ VPWR _1538_ VGND _1464_ _1473_ sg13g2_o21ai_1
XFILLER_49_509 VPWR VGND sg13g2_decap_8
XFILLER_18_907 VPWR VGND sg13g2_decap_8
XFILLER_17_406 VPWR VGND sg13g2_decap_4
XFILLER_45_748 VPWR VGND sg13g2_fill_1
XFILLER_44_225 VPWR VGND sg13g2_fill_1
XFILLER_26_951 VPWR VGND sg13g2_decap_8
XFILLER_13_601 VPWR VGND sg13g2_decap_8
XFILLER_16_52 VPWR VGND sg13g2_fill_1
XFILLER_12_100 VPWR VGND sg13g2_decap_8
XFILLER_41_976 VPWR VGND sg13g2_decap_8
XFILLER_40_431 VPWR VGND sg13g2_fill_1
X_5512__237 VPWR VGND net237 sg13g2_tiehi
XFILLER_10_1020 VPWR VGND sg13g2_decap_8
XFILLER_5_888 VPWR VGND sg13g2_decap_8
XFILLER_35_247 VPWR VGND sg13g2_decap_4
X_3960_ VGND VPWR _2165_ net650 _0199_ _1008_ sg13g2_a21oi_1
XFILLER_17_995 VPWR VGND sg13g2_decap_8
X_2911_ VPWR _2265_ ppwm_i.u_ppwm.global_counter\[12\] VGND sg13g2_inv_1
X_3891_ net835 VPWR _0974_ VGND net522 net669 sg13g2_o21ai_1
XFILLER_32_954 VPWR VGND sg13g2_decap_8
X_2842_ _2196_ net394 VPWR VGND sg13g2_inv_2
X_5561_ net141 VGND VPWR net1138 falu_i.falutop.alu_data_in\[7\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_2
X_5328__45 VPWR VGND net45 sg13g2_tiehi
X_4512_ _1462_ net731 net725 VPWR VGND sg13g2_nand2_1
X_5492_ net297 VGND VPWR _0251_ falu_i.falutop.alu_inst.op\[3\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
Xhold115 falu_i.falutop.div_inst.a\[3\] VPWR VGND net487 sg13g2_dlygate4sd3_1
Xhold104 _0338_ VPWR VGND net476 sg13g2_dlygate4sd3_1
Xhold126 falu_i.falutop.div_inst.acc\[1\] VPWR VGND net498 sg13g2_dlygate4sd3_1
X_5563__124 VPWR VGND net124 sg13g2_tiehi
Xhold159 _0145_ VPWR VGND net531 sg13g2_dlygate4sd3_1
X_4443_ _1395_ _1393_ _1394_ VPWR VGND sg13g2_nand2b_1
Xhold137 _0125_ VPWR VGND net509 sg13g2_dlygate4sd3_1
Xhold148 ppwm_i.u_ppwm.u_pwm.cmp_value\[2\] VPWR VGND net520 sg13g2_dlygate4sd3_1
Xfanout606 _1106_ net606 VPWR VGND sg13g2_buf_8
X_4374_ _1304_ _1321_ _1327_ VPWR VGND sg13g2_nor2_2
X_3325_ VPWR _0068_ _0504_ VGND sg13g2_inv_1
Xfanout639 net640 net639 VPWR VGND sg13g2_buf_1
Xfanout628 net629 net628 VPWR VGND sg13g2_buf_8
Xfanout617 net621 net617 VPWR VGND sg13g2_buf_8
X_3256_ _0445_ _0446_ _0057_ VPWR VGND sg13g2_nor2_1
XFILLER_39_531 VPWR VGND sg13g2_decap_8
XFILLER_39_575 VPWR VGND sg13g2_decap_8
X_3187_ net807 VPWR _0401_ VGND net1111 _0399_ sg13g2_o21ai_1
XFILLER_42_729 VPWR VGND sg13g2_fill_1
XFILLER_35_792 VPWR VGND sg13g2_decap_4
XFILLER_23_954 VPWR VGND sg13g2_decap_8
XFILLER_10_604 VPWR VGND sg13g2_fill_1
X_5567__89 VPWR VGND net89 sg13g2_tiehi
XFILLER_2_869 VPWR VGND sg13g2_decap_8
XFILLER_40_1002 VPWR VGND sg13g2_decap_8
XFILLER_45_523 VPWR VGND sg13g2_fill_1
XFILLER_17_214 VPWR VGND sg13g2_decap_4
XFILLER_26_770 VPWR VGND sg13g2_fill_1
XFILLER_41_740 VPWR VGND sg13g2_fill_2
XFILLER_14_943 VPWR VGND sg13g2_decap_8
XFILLER_4_22 VPWR VGND sg13g2_decap_4
X_3110_ _0350_ _0349_ VPWR VGND falu_i.falutop.i2c_inst.counter\[4\] sg13g2_nand2b_2
X_4090_ net805 VPWR _1094_ VGND net996 _1048_ sg13g2_o21ai_1
XFILLER_49_873 VPWR VGND sg13g2_decap_8
X_3041_ _2395_ net691 _2189_ net694 _2184_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_718 VPWR VGND sg13g2_decap_8
X_4992_ _1899_ VPWR _1934_ VGND _1847_ _1900_ sg13g2_o21ai_1
X_5493__295 VPWR VGND net295 sg13g2_tiehi
XFILLER_23_239 VPWR VGND sg13g2_decap_4
X_3943_ net837 VPWR _1000_ VGND ppwm_i.u_ppwm.u_mem.memory\[91\] net673 sg13g2_o21ai_1
X_5530__145 VPWR VGND net145 sg13g2_tiehi
XFILLER_20_902 VPWR VGND sg13g2_decap_8
XFILLER_32_784 VPWR VGND sg13g2_fill_2
X_3874_ VGND VPWR _2196_ net646 _0156_ _0965_ sg13g2_a21oi_1
X_2825_ VPWR _2179_ net545 VGND sg13g2_inv_1
XFILLER_31_294 VPWR VGND sg13g2_fill_2
Xclkbuf_3_2__f_clk clknet_0_clk clknet_3_2__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_20_979 VPWR VGND sg13g2_decap_8
X_5544_ net363 VGND VPWR net1034 falu_i.falutop.i2c_inst.result\[8\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_5475_ net335 VGND VPWR net851 falu_i.falutop.data_in\[6\] clknet_leaf_5_clk sg13g2_dfrbpq_2
X_4426_ _1220_ _1233_ _1378_ VPWR VGND sg13g2_nor2_1
X_4357_ VPWR _1310_ _1309_ VGND sg13g2_inv_1
X_3308_ _0478_ VPWR _0489_ VGND net700 net696 sg13g2_o21ai_1
X_4288_ _1241_ net714 falu_i.falutop.alu_data_in\[7\] VPWR VGND sg13g2_nand2_2
XFILLER_24_1019 VPWR VGND sg13g2_decap_8
X_3239_ VGND VPWR _2269_ _0433_ _0436_ net795 sg13g2_a21oi_1
XFILLER_39_361 VPWR VGND sg13g2_fill_2
XFILLER_27_534 VPWR VGND sg13g2_decap_8
XFILLER_42_504 VPWR VGND sg13g2_decap_8
XFILLER_42_526 VPWR VGND sg13g2_fill_1
XFILLER_23_751 VPWR VGND sg13g2_decap_8
XFILLER_11_902 VPWR VGND sg13g2_decap_8
XFILLER_13_42 VPWR VGND sg13g2_fill_1
XFILLER_6_427 VPWR VGND sg13g2_fill_2
XFILLER_11_979 VPWR VGND sg13g2_decap_8
XFILLER_2_644 VPWR VGND sg13g2_decap_8
Xhold490 _0314_ VPWR VGND net1142 sg13g2_dlygate4sd3_1
XFILLER_18_534 VPWR VGND sg13g2_decap_8
XFILLER_14_751 VPWR VGND sg13g2_fill_1
XFILLER_14_773 VPWR VGND sg13g2_decap_8
XFILLER_14_795 VPWR VGND sg13g2_decap_8
XFILLER_9_276 VPWR VGND sg13g2_decap_4
X_3590_ _2269_ net592 _0760_ VPWR VGND sg13g2_nor2_1
XFILLER_6_983 VPWR VGND sg13g2_decap_8
X_5260_ net175 VGND VPWR _0022_ falu_i.falutop.i2c_inst.data_in\[18\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_4211_ VGND VPWR net633 _1179_ _0278_ _1180_ sg13g2_a21oi_1
X_5560__149 VPWR VGND net149 sg13g2_tiehi
X_5191_ net1081 falu_i.falutop.data_in\[0\] net624 _0329_ VPWR VGND sg13g2_mux2_1
X_4142_ net525 falu_i.falutop.div_inst.busy _1138_ VPWR VGND sg13g2_and2_1
X_4073_ net861 falu_i.falutop.data_in\[14\] net687 _0242_ VPWR VGND sg13g2_mux2_1
X_3024_ VPWR VGND _2162_ _2377_ net695 _2157_ _2378_ net702 sg13g2_a221oi_1
XFILLER_36_353 VPWR VGND sg13g2_fill_2
X_4975_ _1918_ _1892_ _1917_ VPWR VGND sg13g2_xnor2_1
X_3926_ VGND VPWR _2176_ net650 _0182_ _0991_ sg13g2_a21oi_1
X_3857_ net825 VPWR _0957_ VGND net1008 net658 sg13g2_o21ai_1
XFILLER_20_765 VPWR VGND sg13g2_fill_1
X_2808_ _2162_ net392 VPWR VGND sg13g2_inv_2
X_3788_ VGND VPWR _2225_ net653 _0113_ _0922_ sg13g2_a21oi_1
X_5527_ net165 VGND VPWR net397 falu_i.falutop.div_inst.acc_next\[0\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_5458_ net54 VGND VPWR net1157 ppwm_i.u_ppwm.u_mem.bit_count\[5\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_5389_ net274 VGND VPWR _0148_ ppwm_i.u_ppwm.u_mem.memory\[48\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_2
X_4409_ net616 VPWR _1361_ VGND net767 net566 sg13g2_o21ai_1
XFILLER_39_191 VPWR VGND sg13g2_fill_1
XFILLER_27_331 VPWR VGND sg13g2_fill_1
XFILLER_15_526 VPWR VGND sg13g2_fill_2
XFILLER_27_397 VPWR VGND sg13g2_fill_1
XFILLER_42_356 VPWR VGND sg13g2_fill_1
XFILLER_11_721 VPWR VGND sg13g2_fill_2
XFILLER_11_754 VPWR VGND sg13g2_fill_1
XFILLER_10_286 VPWR VGND sg13g2_fill_1
XFILLER_7_769 VPWR VGND sg13g2_decap_8
XFILLER_3_931 VPWR VGND sg13g2_decap_8
XFILLER_49_71 VPWR VGND sg13g2_decap_4
XFILLER_19_821 VPWR VGND sg13g2_decap_8
XFILLER_46_673 VPWR VGND sg13g2_fill_2
XFILLER_19_898 VPWR VGND sg13g2_decap_8
XFILLER_21_507 VPWR VGND sg13g2_fill_2
XFILLER_33_356 VPWR VGND sg13g2_decap_4
X_4760_ _1707_ _1685_ _1706_ VPWR VGND sg13g2_xnor2_1
X_3711_ net578 VPWR _0871_ VGND ppwm_i.u_ppwm.pwm_value\[6\] net581 sg13g2_o21ai_1
X_4691_ _1563_ VPWR _1639_ VGND _1494_ _1564_ sg13g2_o21ai_1
X_5351__350 VPWR VGND net350 sg13g2_tiehi
X_3642_ _0615_ _0801_ _0805_ _0808_ _0809_ VPWR VGND sg13g2_nor4_1
X_5312_ net77 VGND VPWR _0071_ ppwm_i.u_ppwm.polarity clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3573_ VGND VPWR net578 _0743_ _0744_ net572 sg13g2_a21oi_1
XFILLER_6_780 VPWR VGND sg13g2_fill_1
XFILLER_46_0 VPWR VGND sg13g2_decap_4
X_5243_ net209 VGND VPWR _0005_ falu_i.falutop.i2c_inst.data_in\[1\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_5174_ VGND VPWR _2303_ net617 _0317_ _2104_ sg13g2_a21oi_1
Xhold19 _0191_ VPWR VGND net391 sg13g2_dlygate4sd3_1
X_4125_ _1126_ _1125_ _1112_ _1127_ VPWR VGND sg13g2_a21o_1
XFILLER_29_618 VPWR VGND sg13g2_fill_1
X_4056_ _2294_ _1074_ _1077_ VPWR VGND sg13g2_nor2_1
X_3007_ _2346_ _2360_ _2361_ VPWR VGND sg13g2_nor2_1
XFILLER_37_695 VPWR VGND sg13g2_decap_8
X_4958_ _1901_ _1847_ _1900_ VPWR VGND sg13g2_xnor2_1
X_3909_ net840 VPWR _0983_ VGND ppwm_i.u_ppwm.u_mem.memory\[74\] net678 sg13g2_o21ai_1
X_4889_ VGND VPWR _1832_ _1834_ _1833_ net631 sg13g2_a21oi_2
XFILLER_10_10 VPWR VGND sg13g2_decap_4
X_5508__253 VPWR VGND net253 sg13g2_tiehi
XFILLER_0_967 VPWR VGND sg13g2_decap_8
XFILLER_48_949 VPWR VGND sg13g2_decap_8
XFILLER_15_312 VPWR VGND sg13g2_fill_1
XFILLER_16_846 VPWR VGND sg13g2_decap_8
X_5257__181 VPWR VGND net181 sg13g2_tiehi
XFILLER_7_511 VPWR VGND sg13g2_fill_1
XFILLER_39_905 VPWR VGND sg13g2_fill_2
XFILLER_18_4 VPWR VGND sg13g2_decap_4
XFILLER_47_960 VPWR VGND sg13g2_decap_8
XFILLER_20_1000 VPWR VGND sg13g2_decap_8
X_5379__294 VPWR VGND net294 sg13g2_tiehi
XFILLER_34_676 VPWR VGND sg13g2_fill_1
X_4812_ _1695_ VPWR _1758_ VGND _1693_ _1696_ sg13g2_o21ai_1
XFILLER_22_838 VPWR VGND sg13g2_decap_8
XFILLER_33_164 VPWR VGND sg13g2_decap_8
X_4743_ _1688_ _1529_ _1690_ VPWR VGND sg13g2_xor2_1
X_5566__100 VPWR VGND net100 sg13g2_tiehi
X_4674_ _1622_ net724 net753 VPWR VGND sg13g2_nand2_1
X_3625_ _0792_ VPWR _0793_ VGND _2267_ net591 sg13g2_o21ai_1
X_3556_ net822 VPWR _0728_ VGND net1181 _0614_ sg13g2_o21ai_1
X_5226_ net487 net625 _2135_ VPWR VGND sg13g2_nor2_1
X_3487_ VGND VPWR ppwm_i.u_ppwm.global_counter\[11\] net594 _0662_ _0661_ sg13g2_a21oi_1
X_5157_ falu_i.falutop.data_in\[14\] _1078_ _2093_ _2094_ VPWR VGND sg13g2_nor3_1
XFILLER_29_404 VPWR VGND sg13g2_decap_8
XFILLER_29_437 VPWR VGND sg13g2_fill_2
XFILLER_45_908 VPWR VGND sg13g2_decap_8
XFILLER_38_960 VPWR VGND sg13g2_decap_8
X_4108_ falu_i.falutop.div_inst.acc\[7\] falu_i.falutop.div_inst.b1\[7\] _1110_ VPWR
+ VGND sg13g2_xor2_1
X_5088_ _2028_ net747 net714 falu_i.falutop.alu_data_in\[7\] _2297_ VPWR VGND sg13g2_a22oi_1
XFILLER_44_429 VPWR VGND sg13g2_fill_2
XFILLER_16_109 VPWR VGND sg13g2_fill_1
X_4039_ net816 VPWR _1064_ VGND net1028 _1059_ sg13g2_o21ai_1
XFILLER_13_838 VPWR VGND sg13g2_decap_8
XFILLER_40_668 VPWR VGND sg13g2_fill_2
XFILLER_21_882 VPWR VGND sg13g2_decap_8
XFILLER_20_392 VPWR VGND sg13g2_fill_1
XFILLER_0_720 VPWR VGND sg13g2_decap_4
XFILLER_0_764 VPWR VGND sg13g2_fill_2
XFILLER_47_223 VPWR VGND sg13g2_fill_1
XFILLER_44_930 VPWR VGND sg13g2_decap_8
XFILLER_15_186 VPWR VGND sg13g2_fill_1
XFILLER_12_860 VPWR VGND sg13g2_decap_8
XFILLER_8_853 VPWR VGND sg13g2_decap_8
Xhold308 _0127_ VPWR VGND net960 sg13g2_dlygate4sd3_1
X_3410_ _0584_ _0585_ net591 _0588_ VPWR VGND _0587_ sg13g2_nand4_1
X_4390_ _1342_ VPWR _1343_ VGND net731 _1340_ sg13g2_o21ai_1
Xhold319 ppwm_i.u_ppwm.u_mem.data_sync2 VPWR VGND net971 sg13g2_dlygate4sd3_1
X_3341_ _0519_ _2242_ net784 VPWR VGND sg13g2_nand2_1
X_3272_ VGND VPWR _0457_ _0455_ _2259_ sg13g2_or2_1
X_5011_ _1951_ _1950_ _1953_ VPWR VGND sg13g2_xor2_1
XFILLER_38_245 VPWR VGND sg13g2_fill_2
XFILLER_38_234 VPWR VGND sg13g2_decap_8
XFILLER_19_492 VPWR VGND sg13g2_fill_1
XFILLER_35_963 VPWR VGND sg13g2_decap_8
XFILLER_10_808 VPWR VGND sg13g2_fill_2
X_2987_ _2341_ net692 _2206_ net696 _2215_ VPWR VGND sg13g2_a22oi_1
X_4726_ VGND VPWR _1243_ _1319_ _1673_ _1299_ sg13g2_a21oi_1
X_4657_ _1603_ VPWR _1605_ VGND _1543_ _1545_ sg13g2_o21ai_1
X_3608_ net577 VPWR _0777_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] net590 sg13g2_o21ai_1
X_4588_ _1537_ _1534_ _1535_ VPWR VGND sg13g2_xnor2_1
X_3539_ _0709_ _0710_ _0711_ VPWR VGND sg13g2_nor2b_1
X_5209_ net983 net623 _2123_ VPWR VGND sg13g2_nor2_1
XFILLER_44_204 VPWR VGND sg13g2_fill_1
XFILLER_26_930 VPWR VGND sg13g2_decap_8
X_5551__243 VPWR VGND net243 sg13g2_tiehi
XFILLER_13_613 VPWR VGND sg13g2_fill_1
XFILLER_25_462 VPWR VGND sg13g2_fill_2
XFILLER_41_955 VPWR VGND sg13g2_decap_8
XFILLER_40_454 VPWR VGND sg13g2_decap_8
XFILLER_12_145 VPWR VGND sg13g2_fill_1
XFILLER_16_97 VPWR VGND sg13g2_fill_2
XFILLER_5_867 VPWR VGND sg13g2_decap_8
XFILLER_4_344 VPWR VGND sg13g2_fill_2
XFILLER_35_226 VPWR VGND sg13g2_fill_1
XFILLER_17_974 VPWR VGND sg13g2_decap_8
XFILLER_32_933 VPWR VGND sg13g2_decap_8
X_2910_ VPWR _2264_ ppwm_i.u_ppwm.global_counter\[13\] VGND sg13g2_inv_1
X_3890_ VGND VPWR _2190_ net647 _0164_ _0973_ sg13g2_a21oi_1
X_2841_ VPWR _2195_ net557 VGND sg13g2_inv_1
XFILLER_31_487 VPWR VGND sg13g2_decap_8
X_5560_ net149 VGND VPWR _0319_ falu_i.falutop.alu_data_in\[6\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
XFILLER_8_683 VPWR VGND sg13g2_decap_8
XFILLER_8_650 VPWR VGND sg13g2_fill_1
X_4511_ net760 net730 net566 _1461_ VPWR VGND sg13g2_mux2_1
X_5491_ net299 VGND VPWR _0250_ falu_i.falutop.alu_inst.op\[2\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
XFILLER_7_193 VPWR VGND sg13g2_decap_4
Xhold116 _0339_ VPWR VGND net488 sg13g2_dlygate4sd3_1
X_4442_ VGND VPWR net740 net726 _1394_ net767 sg13g2_a21oi_1
Xhold105 ppwm_i.u_ppwm.u_mem.memory\[22\] VPWR VGND net477 sg13g2_dlygate4sd3_1
Xhold127 _0287_ VPWR VGND net499 sg13g2_dlygate4sd3_1
Xhold149 _0026_ VPWR VGND net521 sg13g2_dlygate4sd3_1
Xhold138 ppwm_i.u_ppwm.u_mem.memory\[85\] VPWR VGND net510 sg13g2_dlygate4sd3_1
X_4373_ _1323_ VPWR _1326_ VGND net744 _1325_ sg13g2_o21ai_1
X_3324_ _0504_ _0502_ _0503_ _0493_ net788 VPWR VGND sg13g2_a22oi_1
Xfanout629 _1076_ net629 VPWR VGND sg13g2_buf_2
Xfanout607 _1105_ net607 VPWR VGND sg13g2_buf_8
Xfanout618 net621 net618 VPWR VGND sg13g2_buf_8
X_3255_ net812 VPWR _0446_ VGND net1134 _0444_ sg13g2_o21ai_1
XFILLER_27_727 VPWR VGND sg13g2_fill_2
X_3186_ net1111 _0399_ _0400_ VPWR VGND sg13g2_and2_1
XFILLER_26_226 VPWR VGND sg13g2_decap_8
XFILLER_27_738 VPWR VGND sg13g2_fill_1
XFILLER_27_749 VPWR VGND sg13g2_fill_1
XFILLER_22_410 VPWR VGND sg13g2_fill_2
XFILLER_23_933 VPWR VGND sg13g2_decap_8
XFILLER_22_454 VPWR VGND sg13g2_fill_1
XFILLER_22_465 VPWR VGND sg13g2_fill_1
XFILLER_10_649 VPWR VGND sg13g2_decap_8
X_4709_ _1655_ _1595_ _1656_ VPWR VGND sg13g2_xor2_1
X_5581__247 VPWR VGND net247 sg13g2_tiehi
XFILLER_2_848 VPWR VGND sg13g2_decap_8
X_5429__176 VPWR VGND net176 sg13g2_tiehi
X_5291__115 VPWR VGND net115 sg13g2_tiehi
X_5436__147 VPWR VGND net147 sg13g2_tiehi
XFILLER_14_922 VPWR VGND sg13g2_decap_8
XFILLER_25_270 VPWR VGND sg13g2_fill_2
XFILLER_14_999 VPWR VGND sg13g2_decap_8
XFILLER_41_796 VPWR VGND sg13g2_fill_1
XFILLER_13_487 VPWR VGND sg13g2_decap_8
X_5443__118 VPWR VGND net118 sg13g2_tiehi
XFILLER_49_852 VPWR VGND sg13g2_decap_8
XFILLER_49_841 VPWR VGND sg13g2_fill_1
XFILLER_49_830 VPWR VGND sg13g2_decap_4
X_3040_ _2392_ _2393_ _2391_ _2394_ VPWR VGND sg13g2_nand3_1
XFILLER_36_579 VPWR VGND sg13g2_fill_1
X_4991_ _1916_ VPWR _1933_ VGND _1892_ _1917_ sg13g2_o21ai_1
XFILLER_16_281 VPWR VGND sg13g2_decap_4
X_3942_ VGND VPWR _2171_ net672 _0190_ _0999_ sg13g2_a21oi_1
XFILLER_17_1016 VPWR VGND sg13g2_decap_8
XFILLER_17_1027 VPWR VGND sg13g2_fill_2
X_3873_ net835 VPWR _0965_ VGND ppwm_i.u_ppwm.u_mem.memory\[57\] net646 sg13g2_o21ai_1
X_2824_ VPWR _2178_ ppwm_i.u_ppwm.u_mem.memory\[80\] VGND sg13g2_inv_1
XFILLER_20_958 VPWR VGND sg13g2_decap_8
XFILLER_31_273 VPWR VGND sg13g2_decap_4
X_5543_ net36 VGND VPWR net1042 falu_i.falutop.i2c_inst.result\[7\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
XFILLER_8_480 VPWR VGND sg13g2_decap_8
X_5474_ net337 VGND VPWR net870 falu_i.falutop.data_in\[5\] clknet_leaf_10_clk sg13g2_dfrbpq_2
X_4425_ _1377_ _1329_ _1332_ _1376_ VPWR VGND sg13g2_and3_1
X_4356_ net772 _2300_ _1304_ _1309_ VPWR VGND sg13g2_nor3_2
X_3307_ VGND VPWR net1162 _0487_ _0488_ _0484_ sg13g2_a21oi_1
X_5361__330 VPWR VGND net330 sg13g2_tiehi
X_4287_ net714 falu_i.falutop.alu_data_in\[7\] _1240_ VPWR VGND sg13g2_nor2_2
X_3238_ _2269_ _0433_ _0435_ VPWR VGND sg13g2_nor2_1
X_3169_ net810 VPWR _0390_ VGND ppwm_i.u_ppwm.pwm_value\[3\] net681 sg13g2_o21ai_1
XFILLER_23_730 VPWR VGND sg13g2_decap_8
XFILLER_11_958 VPWR VGND sg13g2_decap_8
XFILLER_22_295 VPWR VGND sg13g2_fill_2
Xhold480 falu_i.falutop.i2c_inst.counter\[0\] VPWR VGND net1132 sg13g2_dlygate4sd3_1
X_5315__71 VPWR VGND net71 sg13g2_tiehi
XFILLER_49_104 VPWR VGND sg13g2_decap_8
Xhold491 ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] VPWR VGND net1143 sg13g2_dlygate4sd3_1
X_5330__41 VPWR VGND net41 sg13g2_tiehi
XFILLER_1_199 VPWR VGND sg13g2_fill_2
XFILLER_45_321 VPWR VGND sg13g2_fill_1
XFILLER_18_513 VPWR VGND sg13g2_fill_2
XFILLER_18_557 VPWR VGND sg13g2_fill_2
XFILLER_46_888 VPWR VGND sg13g2_decap_8
XFILLER_33_505 VPWR VGND sg13g2_fill_2
XFILLER_14_785 VPWR VGND sg13g2_decap_4
XFILLER_9_244 VPWR VGND sg13g2_decap_8
XFILLER_9_266 VPWR VGND sg13g2_fill_2
XFILLER_6_962 VPWR VGND sg13g2_decap_8
XFILLER_47_1009 VPWR VGND sg13g2_decap_8
XFILLER_5_461 VPWR VGND sg13g2_fill_2
X_4210_ net806 VPWR _1180_ VGND net1100 net633 sg13g2_o21ai_1
X_5190_ net776 net710 net617 _0328_ VPWR VGND sg13g2_mux2_1
X_4141_ _0251_ _2300_ net619 net833 _2292_ VPWR VGND sg13g2_a22oi_1
X_4072_ net894 falu_i.falutop.data_in\[13\] net684 _0241_ VPWR VGND sg13g2_mux2_1
X_3023_ ppwm_i.u_ppwm.u_mem.memory\[89\] net792 net794 _2377_ VPWR VGND sg13g2_nor3_1
XFILLER_36_365 VPWR VGND sg13g2_fill_1
X_4974_ _1917_ _1893_ _1915_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_398 VPWR VGND sg13g2_decap_8
X_3925_ net841 VPWR _0991_ VGND net930 net649 sg13g2_o21ai_1
X_3856_ VGND VPWR _2202_ net642 _0147_ _0956_ sg13g2_a21oi_1
XFILLER_20_744 VPWR VGND sg13g2_decap_8
X_3787_ net824 VPWR _0922_ VGND ppwm_i.u_ppwm.u_mem.memory\[13\] net653 sg13g2_o21ai_1
X_2807_ VPWR _2161_ net914 VGND sg13g2_inv_1
X_5389__274 VPWR VGND net274 sg13g2_tiehi
X_5526_ net169 VGND VPWR _0285_ falu_i.falutop.div_inst.quo\[6\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_5457_ net58 VGND VPWR net1012 ppwm_i.u_ppwm.u_mem.bit_count\[4\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
X_4408_ _1358_ _1359_ _1261_ _1360_ VPWR VGND sg13g2_nand3_1
X_5388_ net276 VGND VPWR _0147_ ppwm_i.u_ppwm.u_mem.memory\[47\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
XFILLER_8_1014 VPWR VGND sg13g2_decap_8
X_4339_ _1292_ _1291_ net710 VPWR VGND sg13g2_nand2b_1
XFILLER_28_822 VPWR VGND sg13g2_fill_1
XFILLER_42_313 VPWR VGND sg13g2_fill_1
XFILLER_10_243 VPWR VGND sg13g2_fill_2
XFILLER_11_744 VPWR VGND sg13g2_fill_2
XFILLER_7_748 VPWR VGND sg13g2_fill_1
XFILLER_6_214 VPWR VGND sg13g2_fill_1
XFILLER_10_265 VPWR VGND sg13g2_fill_1
XFILLER_11_777 VPWR VGND sg13g2_decap_8
XFILLER_11_799 VPWR VGND sg13g2_fill_2
XFILLER_3_910 VPWR VGND sg13g2_decap_8
XFILLER_3_987 VPWR VGND sg13g2_decap_8
XFILLER_38_619 VPWR VGND sg13g2_decap_4
XFILLER_19_800 VPWR VGND sg13g2_fill_1
Xfanout790 net1193 net790 VPWR VGND sg13g2_buf_8
XFILLER_18_354 VPWR VGND sg13g2_fill_2
XFILLER_19_877 VPWR VGND sg13g2_decap_8
XFILLER_45_195 VPWR VGND sg13g2_fill_1
XFILLER_33_324 VPWR VGND sg13g2_fill_1
XFILLER_21_519 VPWR VGND sg13g2_decap_8
X_3710_ VGND VPWR _0870_ _0869_ _0868_ sg13g2_or2_1
XFILLER_41_390 VPWR VGND sg13g2_decap_8
X_4690_ _1638_ _1549_ _1637_ VPWR VGND sg13g2_xnor2_1
X_3641_ VGND VPWR net590 _0806_ _0808_ _0807_ sg13g2_a21oi_1
X_3572_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] _0742_ net588 _0743_ VPWR VGND sg13g2_mux2_1
X_5311_ net79 VGND VPWR _0070_ ppwm_i.u_ppwm.u_ex.cmp_flag_q clknet_leaf_17_clk sg13g2_dfrbpq_2
X_5242_ net211 VGND VPWR _0004_ falu_i.falutop.i2c_inst.data_in\[0\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
XFILLER_39_0 VPWR VGND sg13g2_decap_4
X_5173_ net1114 net617 _2104_ VPWR VGND sg13g2_nor2_1
X_4124_ _1126_ falu_i.falutop.div_inst.b1\[5\] falu_i.falutop.div_inst.acc\[5\] VPWR
+ VGND sg13g2_xnor2_1
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
X_4055_ _1076_ net639 falu_i.falutop.div_inst.done VPWR VGND sg13g2_nand2b_1
X_3006_ _2353_ _2350_ _2359_ _2360_ VPWR VGND sg13g2_a21o_2
XFILLER_25_814 VPWR VGND sg13g2_decap_8
XFILLER_25_869 VPWR VGND sg13g2_decap_8
XFILLER_36_173 VPWR VGND sg13g2_fill_1
X_4957_ _1900_ _1894_ _1898_ VPWR VGND sg13g2_xnor2_1
X_3908_ VGND VPWR _2183_ net678 _0173_ _0982_ sg13g2_a21oi_1
X_4888_ VGND VPWR net632 net565 _1833_ _1276_ sg13g2_a21oi_1
X_3839_ net825 VPWR _0948_ VGND net422 net656 sg13g2_o21ai_1
XFILLER_4_707 VPWR VGND sg13g2_fill_2
X_5509_ net249 VGND VPWR _0268_ falu_i.falutop.div_inst.val\[4\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
XFILLER_0_946 VPWR VGND sg13g2_decap_8
XFILLER_48_928 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_39_clk clknet_3_1__leaf_clk clknet_leaf_39_clk VPWR VGND sg13g2_buf_8
XFILLER_43_611 VPWR VGND sg13g2_decap_8
XFILLER_16_825 VPWR VGND sg13g2_decap_8
X_5454__70 VPWR VGND net70 sg13g2_tiehi
XFILLER_43_655 VPWR VGND sg13g2_fill_2
XFILLER_42_132 VPWR VGND sg13g2_decap_4
X_5515__225 VPWR VGND net225 sg13g2_tiehi
XFILLER_15_346 VPWR VGND sg13g2_fill_2
XFILLER_11_552 VPWR VGND sg13g2_decap_4
XFILLER_7_567 VPWR VGND sg13g2_fill_1
XFILLER_7_534 VPWR VGND sg13g2_decap_4
XFILLER_7_578 VPWR VGND sg13g2_decap_4
XFILLER_38_449 VPWR VGND sg13g2_fill_2
XFILLER_46_493 VPWR VGND sg13g2_decap_4
XFILLER_18_184 VPWR VGND sg13g2_decap_8
X_4811_ _1756_ _1750_ _1757_ VPWR VGND sg13g2_xor2_1
XFILLER_22_817 VPWR VGND sg13g2_decap_8
X_4742_ _1689_ _1688_ _1529_ VPWR VGND sg13g2_nand2b_1
X_4673_ _1621_ net746 net750 VPWR VGND sg13g2_nand2_1
X_3624_ _0792_ ppwm_i.u_ppwm.global_counter\[18\] net591 VPWR VGND sg13g2_nand2_1
X_3555_ net572 _0713_ _0722_ _0726_ _0727_ VPWR VGND sg13g2_nor4_1
X_3486_ net594 ppwm_i.u_ppwm.global_counter\[1\] _0661_ VPWR VGND sg13g2_nor2b_1
X_5225_ _2090_ net776 _2134_ VPWR VGND sg13g2_nor2b_1
X_5156_ _2093_ _2092_ falu_i.falutop.data_in\[13\] VPWR VGND sg13g2_nand2b_1
XFILLER_5_1028 VPWR VGND sg13g2_fill_1
X_5087_ VPWR _2027_ _2026_ VGND sg13g2_inv_1
X_4107_ VGND VPWR net606 _1108_ _0245_ _1109_ sg13g2_a21oi_1
X_4038_ _1050_ _1062_ _1063_ VPWR VGND sg13g2_nor2_1
XFILLER_25_622 VPWR VGND sg13g2_decap_8
XFILLER_24_143 VPWR VGND sg13g2_fill_2
XFILLER_24_154 VPWR VGND sg13g2_fill_1
XFILLER_40_658 VPWR VGND sg13g2_fill_1
XFILLER_21_861 VPWR VGND sg13g2_decap_8
XFILLER_20_371 VPWR VGND sg13g2_fill_1
XFILLER_20_382 VPWR VGND sg13g2_fill_1
XFILLER_21_87 VPWR VGND sg13g2_fill_1
XFILLER_0_710 VPWR VGND sg13g2_fill_2
XFILLER_0_743 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_47_202 VPWR VGND sg13g2_decap_8
XFILLER_35_408 VPWR VGND sg13g2_decap_8
XFILLER_35_419 VPWR VGND sg13g2_fill_1
XFILLER_44_986 VPWR VGND sg13g2_decap_8
XFILLER_16_666 VPWR VGND sg13g2_decap_8
XFILLER_16_677 VPWR VGND sg13g2_fill_1
XFILLER_30_113 VPWR VGND sg13g2_decap_8
XFILLER_30_135 VPWR VGND sg13g2_fill_1
XFILLER_31_647 VPWR VGND sg13g2_fill_2
XFILLER_8_832 VPWR VGND sg13g2_decap_8
XFILLER_8_821 VPWR VGND sg13g2_fill_1
XFILLER_8_810 VPWR VGND sg13g2_decap_8
XFILLER_7_375 VPWR VGND sg13g2_fill_2
Xhold309 ppwm_i.u_ppwm.u_mem.memory\[97\] VPWR VGND net961 sg13g2_dlygate4sd3_1
X_3340_ net782 _2244_ _0518_ VPWR VGND sg13g2_nor2_1
X_3271_ net990 _0456_ _0062_ VPWR VGND sg13g2_nor2_1
X_5010_ _1803_ _1949_ _1951_ _1952_ VPWR VGND sg13g2_nor3_1
XFILLER_39_769 VPWR VGND sg13g2_fill_2
XFILLER_38_268 VPWR VGND sg13g2_decap_8
X_5496__283 VPWR VGND net283 sg13g2_tiehi
XFILLER_21_179 VPWR VGND sg13g2_decap_4
X_2986_ VPWR VGND _2225_ _2338_ net693 _2220_ _2340_ net704 sg13g2_a221oi_1
X_4725_ VGND VPWR _1244_ _1383_ _1672_ _1313_ sg13g2_a21oi_1
X_4656_ _1543_ _1545_ _1603_ _1604_ VPWR VGND sg13g2_nor3_1
X_3607_ VGND VPWR ppwm_i.u_ppwm.global_counter\[17\] net591 _0776_ _0775_ sg13g2_a21oi_1
X_4587_ _1536_ _1534_ _1535_ VPWR VGND sg13g2_nand2b_1
XFILLER_1_507 VPWR VGND sg13g2_decap_8
X_3538_ VGND VPWR _0688_ _0690_ _0710_ _0689_ sg13g2_a21oi_1
X_3469_ net573 _0638_ _0642_ _0644_ _0645_ VPWR VGND sg13g2_nor4_1
X_5208_ _2098_ net777 _2122_ VPWR VGND sg13g2_nor2b_1
X_5139_ _2027_ VPWR _2077_ VGND _2025_ _2056_ sg13g2_o21ai_1
XFILLER_17_419 VPWR VGND sg13g2_decap_8
XFILLER_38_780 VPWR VGND sg13g2_decap_8
X_5371__310 VPWR VGND net310 sg13g2_tiehi
XFILLER_41_934 VPWR VGND sg13g2_decap_8
XFILLER_26_986 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_fill_1
XFILLER_32_20 VPWR VGND sg13g2_fill_1
XFILLER_40_499 VPWR VGND sg13g2_decap_8
XFILLER_40_488 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_fill_2
XFILLER_5_846 VPWR VGND sg13g2_decap_8
XFILLER_48_555 VPWR VGND sg13g2_decap_4
XFILLER_35_205 VPWR VGND sg13g2_fill_1
XFILLER_17_953 VPWR VGND sg13g2_decap_8
XFILLER_44_783 VPWR VGND sg13g2_decap_4
XFILLER_31_411 VPWR VGND sg13g2_decap_8
X_2840_ VPWR _2194_ net866 VGND sg13g2_inv_1
XFILLER_32_989 VPWR VGND sg13g2_decap_8
X_4510_ VPWR VGND _1460_ _1457_ _1459_ _1412_ _0297_ _1456_ sg13g2_a221oi_1
X_5490_ net301 VGND VPWR _0249_ falu_i.falutop.alu_inst.op\[1\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_2
Xhold117 falu_i.falutop.div_inst.acc\[2\] VPWR VGND net489 sg13g2_dlygate4sd3_1
X_4441_ _1393_ net726 _1232_ VPWR VGND sg13g2_nand2_2
Xhold106 _0121_ VPWR VGND net478 sg13g2_dlygate4sd3_1
Xhold128 ppwm_i.u_ppwm.u_mem.memory\[101\] VPWR VGND net500 sg13g2_dlygate4sd3_1
Xhold139 _0185_ VPWR VGND net511 sg13g2_dlygate4sd3_1
X_4372_ VGND VPWR _1325_ _1321_ _1279_ sg13g2_or2_1
X_5348__356 VPWR VGND net356 sg13g2_tiehi
Xfanout608 _2418_ net608 VPWR VGND sg13g2_buf_8
X_3323_ VPWR VGND _0482_ _2422_ _0499_ _0478_ _0503_ _0495_ sg13g2_a221oi_1
Xfanout619 net621 net619 VPWR VGND sg13g2_buf_8
X_3254_ net1134 _0444_ _0445_ VPWR VGND sg13g2_and2_1
XFILLER_2_1009 VPWR VGND sg13g2_decap_8
X_3185_ ppwm_i.u_ppwm.u_mem.bit_count\[3\] ppwm_i.u_ppwm.u_mem.bit_count\[1\] net378
+ _0398_ _0399_ VPWR VGND sg13g2_nor4_1
XFILLER_23_912 VPWR VGND sg13g2_decap_8
XFILLER_23_989 VPWR VGND sg13g2_decap_8
X_2969_ VPWR VGND _2229_ net789 net689 _2234_ _2323_ net698 sg13g2_a221oi_1
X_4708_ _1654_ VPWR _1655_ VGND net749 _1592_ sg13g2_o21ai_1
X_5546__313 VPWR VGND net313 sg13g2_tiehi
X_4639_ _1406_ _1587_ _1588_ VPWR VGND sg13g2_nor2_1
XFILLER_2_827 VPWR VGND sg13g2_decap_8
X_5399__254 VPWR VGND net254 sg13g2_tiehi
XFILLER_14_901 VPWR VGND sg13g2_decap_8
XFILLER_41_742 VPWR VGND sg13g2_fill_1
XFILLER_13_422 VPWR VGND sg13g2_decap_4
XFILLER_41_753 VPWR VGND sg13g2_decap_4
XFILLER_40_241 VPWR VGND sg13g2_fill_2
XFILLER_9_404 VPWR VGND sg13g2_fill_2
XFILLER_13_466 VPWR VGND sg13g2_decap_8
XFILLER_14_978 VPWR VGND sg13g2_decap_8
XFILLER_9_448 VPWR VGND sg13g2_decap_4
XFILLER_5_621 VPWR VGND sg13g2_fill_1
XFILLER_4_186 VPWR VGND sg13g2_fill_2
XFILLER_0_370 VPWR VGND sg13g2_decap_8
XFILLER_1_882 VPWR VGND sg13g2_decap_8
X_4990_ _1931_ _1932_ _0305_ VPWR VGND sg13g2_nor2_1
XFILLER_23_208 VPWR VGND sg13g2_decap_8
XFILLER_23_219 VPWR VGND sg13g2_fill_2
XFILLER_44_580 VPWR VGND sg13g2_fill_1
X_3941_ net838 VPWR _0999_ VGND ppwm_i.u_ppwm.u_mem.memory\[90\] net672 sg13g2_o21ai_1
X_3872_ VGND VPWR _2196_ net671 _0155_ _0964_ sg13g2_a21oi_1
XFILLER_31_241 VPWR VGND sg13g2_fill_2
X_2823_ VPWR _2177_ net948 VGND sg13g2_inv_1
XFILLER_20_937 VPWR VGND sg13g2_decap_8
XFILLER_31_285 VPWR VGND sg13g2_decap_4
XFILLER_32_797 VPWR VGND sg13g2_fill_2
X_5542_ net44 VGND VPWR _0301_ falu_i.falutop.i2c_inst.result\[6\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_31_296 VPWR VGND sg13g2_fill_1
XFILLER_9_993 VPWR VGND sg13g2_decap_8
X_5473_ net339 VGND VPWR net882 falu_i.falutop.data_in\[4\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4424_ _1285_ VPWR _1376_ VGND _1284_ _1286_ sg13g2_o21ai_1
X_4355_ _1308_ net726 _1219_ VPWR VGND sg13g2_nand2_1
X_3306_ _0487_ _0476_ _0485_ VPWR VGND sg13g2_xnor2_1
X_4286_ _1237_ _1238_ _1239_ VPWR VGND sg13g2_and2_1
X_3237_ net1146 _0433_ _0050_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_363 VPWR VGND sg13g2_fill_1
X_3168_ VGND VPWR _2286_ net681 _0026_ _0389_ sg13g2_a21oi_1
XFILLER_14_219 VPWR VGND sg13g2_decap_4
X_3099_ net816 VPWR _2448_ VGND net901 net1002 sg13g2_o21ai_1
XFILLER_11_937 VPWR VGND sg13g2_decap_8
XFILLER_23_786 VPWR VGND sg13g2_decap_8
XFILLER_10_436 VPWR VGND sg13g2_decap_8
XFILLER_6_429 VPWR VGND sg13g2_fill_1
XFILLER_2_635 VPWR VGND sg13g2_decap_4
Xhold481 falu_i.falutop.div_inst.val\[0\] VPWR VGND net1133 sg13g2_dlygate4sd3_1
Xhold470 falu_i.falutop.data_in\[10\] VPWR VGND net1122 sg13g2_dlygate4sd3_1
Xhold492 ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] VPWR VGND net1144 sg13g2_dlygate4sd3_1
XFILLER_38_63 VPWR VGND sg13g2_fill_2
XFILLER_45_300 VPWR VGND sg13g2_decap_8
XFILLER_45_388 VPWR VGND sg13g2_fill_2
XFILLER_45_377 VPWR VGND sg13g2_fill_1
XFILLER_41_583 VPWR VGND sg13g2_fill_1
XFILLER_9_212 VPWR VGND sg13g2_fill_2
XFILLER_13_296 VPWR VGND sg13g2_decap_8
XFILLER_6_941 VPWR VGND sg13g2_decap_8
XFILLER_10_992 VPWR VGND sg13g2_decap_8
X_5267__162 VPWR VGND net162 sg13g2_tiehi
XFILLER_5_495 VPWR VGND sg13g2_fill_2
X_4140_ _0250_ _2299_ net619 net833 _2293_ VPWR VGND sg13g2_a22oi_1
X_4071_ net926 falu_i.falutop.data_in\[12\] net685 _0240_ VPWR VGND sg13g2_mux2_1
XFILLER_23_1010 VPWR VGND sg13g2_decap_8
XFILLER_49_683 VPWR VGND sg13g2_decap_8
X_3022_ VGND VPWR _2167_ net690 _2376_ net709 sg13g2_a21oi_1
XFILLER_36_333 VPWR VGND sg13g2_fill_2
XFILLER_24_528 VPWR VGND sg13g2_decap_4
X_4973_ _1916_ _1893_ _1915_ VPWR VGND sg13g2_nand2_1
XFILLER_17_580 VPWR VGND sg13g2_fill_1
XFILLER_17_591 VPWR VGND sg13g2_fill_2
X_3924_ VGND VPWR _2176_ net677 _0181_ _0990_ sg13g2_a21oi_1
X_3855_ net825 VPWR _0956_ VGND net1008 net642 sg13g2_o21ai_1
X_3786_ VGND VPWR _2226_ net641 _0112_ _0921_ sg13g2_a21oi_1
X_2806_ VPWR _2160_ net528 VGND sg13g2_inv_1
XFILLER_30_1014 VPWR VGND sg13g2_decap_8
X_5525_ net174 VGND VPWR net433 falu_i.falutop.div_inst.quo\[5\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_5456_ net62 VGND VPWR _0215_ ppwm_i.u_ppwm.u_mem.bit_count\[3\] clknet_leaf_4_clk
+ sg13g2_dfrbpq_2
X_4407_ _1359_ _1258_ _1357_ VPWR VGND sg13g2_nand2_1
X_5387_ net278 VGND VPWR _0146_ ppwm_i.u_ppwm.u_mem.memory\[46\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_4338_ _1289_ VPWR _1291_ VGND net730 _1290_ sg13g2_o21ai_1
X_4269_ _1219_ _1221_ _1222_ VPWR VGND sg13g2_nor2_1
XFILLER_27_366 VPWR VGND sg13g2_decap_4
XFILLER_28_878 VPWR VGND sg13g2_decap_4
XFILLER_15_528 VPWR VGND sg13g2_fill_1
XFILLER_23_594 VPWR VGND sg13g2_decap_8
XFILLER_10_255 VPWR VGND sg13g2_fill_1
XFILLER_46_1021 VPWR VGND sg13g2_decap_8
XFILLER_3_966 VPWR VGND sg13g2_decap_8
XFILLER_2_465 VPWR VGND sg13g2_decap_4
XFILLER_1_14 VPWR VGND sg13g2_decap_8
Xfanout780 net887 net780 VPWR VGND sg13g2_buf_2
Xfanout791 net1168 net791 VPWR VGND sg13g2_buf_8
XFILLER_19_856 VPWR VGND sg13g2_decap_8
XFILLER_33_303 VPWR VGND sg13g2_fill_1
XFILLER_34_837 VPWR VGND sg13g2_decap_8
XFILLER_21_509 VPWR VGND sg13g2_fill_1
X_3640_ net579 VPWR _0807_ VGND net1160 net589 sg13g2_o21ai_1
X_3571_ VGND VPWR _2262_ net593 _0742_ _0741_ sg13g2_a21oi_1
X_5310_ net81 VGND VPWR _0069_ ppwm_i.u_ppwm.pc\[3\] clknet_leaf_22_clk sg13g2_dfrbpq_1
XFILLER_5_270 VPWR VGND sg13g2_decap_4
X_5241_ net93 VGND VPWR _0003_ falu_i.falutop.i2c_inst.data_in\[19\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_1
X_5172_ net1135 net760 net618 _0316_ VPWR VGND sg13g2_mux2_1
X_4123_ _1124_ _1123_ _1113_ _1125_ VPWR VGND sg13g2_a21o_1
X_4054_ net380 _1074_ _1075_ VPWR VGND sg13g2_nor2_2
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
X_3005_ VPWR VGND _2358_ net787 _2357_ _2355_ _2359_ _2356_ sg13g2_a221oi_1
XFILLER_25_848 VPWR VGND sg13g2_decap_8
XFILLER_40_818 VPWR VGND sg13g2_decap_8
X_4956_ _1899_ _1894_ _1898_ VPWR VGND sg13g2_nand2_1
XFILLER_33_881 VPWR VGND sg13g2_decap_4
X_3907_ net839 VPWR _0982_ VGND ppwm_i.u_ppwm.u_mem.memory\[73\] net678 sg13g2_o21ai_1
X_4887_ _1240_ _1727_ _1832_ VPWR VGND sg13g2_nor2_1
XFILLER_20_531 VPWR VGND sg13g2_fill_1
X_3838_ VGND VPWR _2208_ net656 _0138_ _0947_ sg13g2_a21oi_1
XFILLER_20_564 VPWR VGND sg13g2_fill_1
X_5508_ net253 VGND VPWR _0267_ falu_i.falutop.div_inst.val\[3\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_3769_ net824 VPWR _0913_ VGND net847 net642 sg13g2_o21ai_1
X_5547__293 VPWR VGND net293 sg13g2_tiehi
X_5439_ net135 VGND VPWR _0198_ ppwm_i.u_ppwm.u_mem.memory\[98\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
XFILLER_0_925 VPWR VGND sg13g2_decap_8
XFILLER_48_907 VPWR VGND sg13g2_decap_8
XFILLER_16_804 VPWR VGND sg13g2_decap_8
XFILLER_42_100 VPWR VGND sg13g2_decap_4
XFILLER_11_586 VPWR VGND sg13g2_fill_1
XFILLER_13_1020 VPWR VGND sg13g2_decap_8
XFILLER_3_796 VPWR VGND sg13g2_decap_8
XFILLER_47_995 VPWR VGND sg13g2_decap_8
X_4810_ VGND VPWR _1688_ _1751_ _1756_ _1755_ sg13g2_a21oi_1
XFILLER_18_196 VPWR VGND sg13g2_decap_8
X_4741_ net719 net769 _1688_ VPWR VGND sg13g2_and2_1
X_4672_ _1561_ _1552_ _1559_ _1620_ VPWR VGND sg13g2_a21o_1
X_3623_ _0757_ _0628_ _0790_ _0791_ VPWR VGND sg13g2_a21o_1
X_3554_ VGND VPWR net588 _0724_ _0726_ _0725_ sg13g2_a21oi_1
X_3485_ VGND VPWR _0619_ _0658_ _0660_ _0659_ sg13g2_a21oi_1
X_5224_ VGND VPWR net625 _2133_ _0338_ _2131_ sg13g2_a21oi_1
X_5155_ falu_i.falutop.data_in\[12\] _2091_ _2092_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_1007 VPWR VGND sg13g2_decap_8
X_5086_ _1241_ _1729_ _2026_ VPWR VGND sg13g2_nor2b_2
X_4106_ net1009 net606 _1109_ VPWR VGND sg13g2_nor2_1
XFILLER_29_439 VPWR VGND sg13g2_fill_1
X_4037_ _2445_ _0343_ _1049_ _1062_ VPWR VGND sg13g2_nor3_1
XFILLER_38_995 VPWR VGND sg13g2_decap_8
XFILLER_37_494 VPWR VGND sg13g2_fill_1
X_5358__336 VPWR VGND net336 sg13g2_tiehi
X_4939_ VGND VPWR _2304_ net563 _1883_ _1282_ sg13g2_a21oi_1
XFILLER_21_840 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_21_22 VPWR VGND sg13g2_decap_8
XFILLER_43_1024 VPWR VGND sg13g2_decap_4
XFILLER_0_733 VPWR VGND sg13g2_fill_2
XFILLER_0_799 VPWR VGND sg13g2_decap_8
XFILLER_29_984 VPWR VGND sg13g2_decap_8
XFILLER_16_623 VPWR VGND sg13g2_decap_8
X_5439__135 VPWR VGND net135 sg13g2_tiehi
XFILLER_44_965 VPWR VGND sg13g2_decap_8
XFILLER_11_350 VPWR VGND sg13g2_fill_1
XFILLER_7_310 VPWR VGND sg13g2_decap_4
XFILLER_7_46 VPWR VGND sg13g2_fill_2
XFILLER_12_895 VPWR VGND sg13g2_decap_8
XFILLER_8_888 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_decap_8
X_5446__106 VPWR VGND net106 sg13g2_tiehi
X_3270_ _0456_ net812 _0455_ VPWR VGND sg13g2_nand2_1
XFILLER_3_571 VPWR VGND sg13g2_decap_8
XFILLER_47_792 VPWR VGND sg13g2_decap_4
XFILLER_35_910 VPWR VGND sg13g2_fill_2
XFILLER_34_486 VPWR VGND sg13g2_decap_8
XFILLER_35_998 VPWR VGND sg13g2_decap_8
X_2985_ VGND VPWR _2230_ net688 _2339_ net788 sg13g2_a21oi_1
X_4724_ _1323_ VPWR _1671_ VGND net748 _1325_ sg13g2_o21ai_1
XFILLER_30_670 VPWR VGND sg13g2_fill_1
X_4655_ _1603_ _1600_ _1601_ VPWR VGND sg13g2_xnor2_1
X_3606_ _2268_ net592 _0775_ VPWR VGND sg13g2_nor2_1
X_4586_ VGND VPWR net721 _1467_ _1535_ _1470_ sg13g2_a21oi_1
X_3537_ _0709_ _2248_ net600 VPWR VGND sg13g2_xnor2_1
XFILLER_27_1008 VPWR VGND sg13g2_decap_8
X_3468_ _0618_ _0643_ _0644_ VPWR VGND sg13g2_nor2_1
X_3399_ VPWR VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] _0576_ _2263_ ppwm_i.u_ppwm.u_ex.reg_value_q\[5\]
+ _0577_ _2262_ sg13g2_a221oi_1
X_5207_ VGND VPWR net623 _2121_ _0333_ _2119_ sg13g2_a21oi_1
X_5138_ VGND VPWR _2055_ _2060_ _2076_ _2062_ sg13g2_a21oi_1
XFILLER_29_236 VPWR VGND sg13g2_decap_4
XFILLER_45_707 VPWR VGND sg13g2_decap_4
X_5069_ _1317_ _2008_ _2010_ VPWR VGND _2009_ sg13g2_nand3b_1
XFILLER_16_11 VPWR VGND sg13g2_decap_8
X_5475__335 VPWR VGND net335 sg13g2_tiehi
XFILLER_26_965 VPWR VGND sg13g2_decap_8
XFILLER_40_401 VPWR VGND sg13g2_fill_1
XFILLER_16_77 VPWR VGND sg13g2_fill_2
XFILLER_25_464 VPWR VGND sg13g2_fill_1
XFILLER_40_423 VPWR VGND sg13g2_fill_2
XFILLER_12_114 VPWR VGND sg13g2_fill_2
XFILLER_13_659 VPWR VGND sg13g2_fill_2
XFILLER_20_191 VPWR VGND sg13g2_fill_2
XFILLER_5_825 VPWR VGND sg13g2_decap_8
XFILLER_4_302 VPWR VGND sg13g2_decap_4
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_36_718 VPWR VGND sg13g2_decap_8
XFILLER_17_932 VPWR VGND sg13g2_decap_8
XFILLER_43_250 VPWR VGND sg13g2_decap_4
XFILLER_16_453 VPWR VGND sg13g2_decap_8
XFILLER_16_464 VPWR VGND sg13g2_fill_1
XFILLER_31_401 VPWR VGND sg13g2_fill_1
XFILLER_32_968 VPWR VGND sg13g2_decap_8
XFILLER_8_630 VPWR VGND sg13g2_decap_4
Xhold107 falu_i.falutop.div_inst.b1\[0\] VPWR VGND net479 sg13g2_dlygate4sd3_1
X_4440_ _1392_ net728 net766 VPWR VGND sg13g2_nand2_1
Xhold118 _0288_ VPWR VGND net490 sg13g2_dlygate4sd3_1
Xhold129 _0200_ VPWR VGND net501 sg13g2_dlygate4sd3_1
XFILLER_4_880 VPWR VGND sg13g2_decap_8
X_4371_ _1279_ _1321_ _1324_ VPWR VGND sg13g2_nor2_2
Xfanout609 net610 net609 VPWR VGND sg13g2_buf_8
X_3322_ _0501_ VPWR _0502_ VGND _2253_ _0499_ sg13g2_o21ai_1
X_3253_ net795 net955 _0444_ _0056_ VPWR VGND sg13g2_nor3_1
XFILLER_39_523 VPWR VGND sg13g2_decap_4
X_3184_ ppwm_i.u_ppwm.u_mem.bit_count\[5\] net1010 net512 _0398_ VPWR VGND _2155_
+ sg13g2_nand4_1
XFILLER_27_729 VPWR VGND sg13g2_fill_1
X_5277__142 VPWR VGND net142 sg13g2_tiehi
XFILLER_35_751 VPWR VGND sg13g2_fill_2
XFILLER_22_412 VPWR VGND sg13g2_fill_1
XFILLER_10_618 VPWR VGND sg13g2_decap_8
XFILLER_23_968 VPWR VGND sg13g2_decap_8
X_2968_ _2322_ net693 _2224_ net701 _2219_ VPWR VGND sg13g2_a22oi_1
XFILLER_33_1023 VPWR VGND sg13g2_decap_4
X_4707_ VGND VPWR _1654_ _1653_ _1652_ sg13g2_or2_1
X_2899_ _2253_ net1162 VPWR VGND sg13g2_inv_2
X_4638_ _1585_ _1586_ _1587_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_806 VPWR VGND sg13g2_decap_8
X_4569_ _1498_ _1503_ _1481_ _1519_ VPWR VGND _1518_ sg13g2_nand4_1
XFILLER_49_309 VPWR VGND sg13g2_decap_4
XFILLER_40_1027 VPWR VGND sg13g2_fill_2
XFILLER_40_1016 VPWR VGND sg13g2_decap_8
XFILLER_26_751 VPWR VGND sg13g2_fill_2
XFILLER_14_957 VPWR VGND sg13g2_decap_8
XFILLER_25_272 VPWR VGND sg13g2_fill_1
XFILLER_43_64 VPWR VGND sg13g2_decap_8
XFILLER_9_427 VPWR VGND sg13g2_decap_8
XFILLER_4_110 VPWR VGND sg13g2_decap_4
XFILLER_5_699 VPWR VGND sg13g2_decap_8
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_49_887 VPWR VGND sg13g2_decap_8
XFILLER_17_773 VPWR VGND sg13g2_fill_2
X_3940_ VGND VPWR _2172_ net646 _0189_ _0998_ sg13g2_a21oi_1
XFILLER_17_795 VPWR VGND sg13g2_decap_4
X_3871_ net835 VPWR _0964_ VGND net398 net665 sg13g2_o21ai_1
XFILLER_20_916 VPWR VGND sg13g2_decap_8
X_2822_ _2176_ net417 VPWR VGND sg13g2_inv_2
X_5541_ net52 VGND VPWR _0300_ falu_i.falutop.i2c_inst.result\[5\] clknet_leaf_40_clk
+ sg13g2_dfrbpq_1
XFILLER_9_972 VPWR VGND sg13g2_decap_8
XFILLER_8_493 VPWR VGND sg13g2_fill_1
X_5472_ net341 VGND VPWR net993 falu_i.falutop.data_in\[3\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4423_ _1375_ _1219_ _1235_ VPWR VGND sg13g2_xnor2_1
X_4354_ _1220_ VPWR _1307_ VGND _1303_ net631 sg13g2_o21ai_1
X_3305_ _0476_ _0485_ _0486_ VPWR VGND sg13g2_nor2_1
X_4285_ VGND VPWR _1238_ net754 net729 sg13g2_or2_1
X_3236_ net813 VPWR _0434_ VGND net1145 _0431_ sg13g2_o21ai_1
X_3167_ net808 VPWR _0389_ VGND ppwm_i.u_ppwm.pwm_value\[2\] net681 sg13g2_o21ai_1
X_3098_ _2437_ _2446_ _2447_ VPWR VGND sg13g2_nor2_1
XFILLER_27_559 VPWR VGND sg13g2_decap_8
XFILLER_11_916 VPWR VGND sg13g2_decap_8
XFILLER_23_765 VPWR VGND sg13g2_decap_8
XFILLER_7_909 VPWR VGND sg13g2_decap_8
XFILLER_22_297 VPWR VGND sg13g2_fill_1
Xhold471 falu_i.falutop.data_in\[9\] VPWR VGND net1123 sg13g2_dlygate4sd3_1
Xhold460 _0401_ VPWR VGND net1112 sg13g2_dlygate4sd3_1
Xhold493 ppwm_i.u_ppwm.global_counter\[5\] VPWR VGND net1145 sg13g2_dlygate4sd3_1
XFILLER_1_135 VPWR VGND sg13g2_fill_1
Xhold482 ppwm_i.u_ppwm.global_counter\[12\] VPWR VGND net1134 sg13g2_dlygate4sd3_1
X_5518__213 VPWR VGND net213 sg13g2_tiehi
XFILLER_18_548 VPWR VGND sg13g2_decap_4
XFILLER_33_507 VPWR VGND sg13g2_fill_1
XFILLER_14_721 VPWR VGND sg13g2_fill_2
XFILLER_13_242 VPWR VGND sg13g2_fill_1
XFILLER_6_920 VPWR VGND sg13g2_decap_8
XFILLER_10_971 VPWR VGND sg13g2_decap_8
XFILLER_6_997 VPWR VGND sg13g2_decap_8
XFILLER_5_463 VPWR VGND sg13g2_fill_1
XFILLER_1_691 VPWR VGND sg13g2_decap_8
X_4070_ net858 falu_i.falutop.data_in\[11\] net685 _0239_ VPWR VGND sg13g2_mux2_1
X_3021_ _2375_ net602 VPWR VGND sg13g2_inv_2
XFILLER_37_824 VPWR VGND sg13g2_decap_8
X_4972_ _1914_ _1901_ _1915_ VPWR VGND sg13g2_xor2_1
X_3923_ net840 VPWR _0990_ VGND ppwm_i.u_ppwm.u_mem.memory\[81\] net677 sg13g2_o21ai_1
X_3854_ VGND VPWR _2202_ net658 _0146_ _0955_ sg13g2_a21oi_1
X_2805_ VPWR _2159_ net445 VGND sg13g2_inv_1
X_3785_ net832 VPWR _0921_ VGND net933 net641 sg13g2_o21ai_1
X_5524_ net178 VGND VPWR net406 falu_i.falutop.div_inst.quo\[4\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_5455_ net66 VGND VPWR net1053 ppwm_i.u_ppwm.u_mem.bit_count\[2\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_4406_ VGND VPWR _1358_ _1357_ _1258_ sg13g2_or2_1
X_5246__203 VPWR VGND net203 sg13g2_tiehi
X_5386_ net280 VGND VPWR net531 ppwm_i.u_ppwm.u_mem.memory\[45\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4337_ net707 net735 _1290_ VPWR VGND sg13g2_nor2_1
X_4268_ net744 net770 _1221_ VPWR VGND sg13g2_nor2_1
X_3219_ net864 _0411_ _0421_ _0422_ _0044_ VPWR VGND sg13g2_nor4_1
XFILLER_28_813 VPWR VGND sg13g2_fill_2
X_4199_ _1170_ VPWR _1171_ VGND net856 net567 sg13g2_o21ai_1
X_5368__316 VPWR VGND net316 sg13g2_tiehi
XFILLER_40_76 VPWR VGND sg13g2_fill_2
XFILLER_46_1000 VPWR VGND sg13g2_decap_8
XFILLER_3_945 VPWR VGND sg13g2_decap_8
XFILLER_2_400 VPWR VGND sg13g2_fill_1
Xhold290 ppwm_i.u_ppwm.global_counter\[1\] VPWR VGND net942 sg13g2_dlygate4sd3_1
Xfanout781 falu_i.falutop.div_inst.start net781 VPWR VGND sg13g2_buf_1
Xfanout770 falu_i.falutop.alu_data_in\[0\] net770 VPWR VGND sg13g2_buf_8
Xfanout792 ppwm_i.u_ppwm.pc\[1\] net792 VPWR VGND sg13g2_buf_8
XFILLER_19_835 VPWR VGND sg13g2_decap_8
XFILLER_46_698 VPWR VGND sg13g2_fill_1
XFILLER_45_186 VPWR VGND sg13g2_fill_2
X_3570_ ppwm_i.u_ppwm.global_counter\[5\] net593 _0741_ VPWR VGND sg13g2_nor2_1
XFILLER_10_790 VPWR VGND sg13g2_decap_8
XFILLER_6_750 VPWR VGND sg13g2_fill_2
X_5240_ VGND VPWR net625 _2145_ _0342_ _2143_ sg13g2_a21oi_1
X_5171_ net1127 net765 net618 _0315_ VPWR VGND sg13g2_mux2_1
X_4122_ _1124_ falu_i.falutop.div_inst.b1\[4\] falu_i.falutop.div_inst.acc\[4\] VPWR
+ VGND sg13g2_xnor2_1
X_5425__192 VPWR VGND net192 sg13g2_tiehi
X_4053_ _2291_ falu_i.falutop.i2c_inst.op\[1\] _2292_ _2293_ _1074_ VPWR VGND sg13g2_or4_1
X_3004_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[44\] net708 net692 ppwm_i.u_ppwm.u_mem.memory\[51\]
+ _2358_ net701 sg13g2_a221oi_1
Xinput3 ui_in[3] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_665 VPWR VGND sg13g2_decap_8
XFILLER_24_315 VPWR VGND sg13g2_fill_1
X_4955_ _1898_ _1895_ _1896_ VPWR VGND sg13g2_xnor2_1
X_3906_ VGND VPWR _2184_ net670 _0172_ _0981_ sg13g2_a21oi_1
X_4886_ _1831_ _1829_ VPWR VGND _1830_ sg13g2_nand2b_2
XFILLER_20_521 VPWR VGND sg13g2_fill_2
X_3837_ net829 VPWR _0947_ VGND ppwm_i.u_ppwm.u_mem.memory\[38\] net656 sg13g2_o21ai_1
X_5432__163 VPWR VGND net163 sg13g2_tiehi
XFILLER_20_598 VPWR VGND sg13g2_decap_8
X_3768_ VGND VPWR _2232_ net659 _0103_ _0912_ sg13g2_a21oi_1
X_5507_ net257 VGND VPWR net979 falu_i.falutop.div_inst.val\[2\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_2
X_3699_ _0859_ VPWR _0860_ VGND _0857_ _0858_ sg13g2_o21ai_1
XFILLER_0_904 VPWR VGND sg13g2_decap_8
X_5438_ net139 VGND VPWR _0197_ ppwm_i.u_ppwm.u_mem.memory\[97\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
X_5369_ net314 VGND VPWR _0128_ ppwm_i.u_ppwm.u_mem.memory\[28\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_47_418 VPWR VGND sg13g2_fill_1
XFILLER_28_621 VPWR VGND sg13g2_fill_1
XFILLER_27_153 VPWR VGND sg13g2_decap_4
XFILLER_43_635 VPWR VGND sg13g2_fill_2
XFILLER_43_624 VPWR VGND sg13g2_decap_8
XFILLER_27_186 VPWR VGND sg13g2_decap_8
XFILLER_35_43 VPWR VGND sg13g2_fill_2
XFILLER_43_657 VPWR VGND sg13g2_fill_1
XFILLER_31_808 VPWR VGND sg13g2_fill_2
XFILLER_24_893 VPWR VGND sg13g2_decap_8
X_5485__315 VPWR VGND net315 sg13g2_tiehi
XFILLER_3_742 VPWR VGND sg13g2_decap_8
XFILLER_2_285 VPWR VGND sg13g2_decap_4
XFILLER_47_974 VPWR VGND sg13g2_decap_8
XFILLER_19_643 VPWR VGND sg13g2_decap_8
XFILLER_20_1014 VPWR VGND sg13g2_decap_8
XFILLER_33_134 VPWR VGND sg13g2_fill_2
XFILLER_33_145 VPWR VGND sg13g2_fill_2
XFILLER_15_882 VPWR VGND sg13g2_decap_8
X_4740_ _1687_ net742 net751 VPWR VGND sg13g2_nand2_1
X_4671_ _1618_ VPWR _1619_ VGND _1374_ _1612_ sg13g2_o21ai_1
X_3622_ net574 _0787_ _0788_ _0789_ _0790_ VPWR VGND sg13g2_nor4_1
X_3553_ net577 VPWR _0725_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] net588 sg13g2_o21ai_1
XFILLER_44_0 VPWR VGND sg13g2_fill_2
X_3484_ net576 VPWR _0659_ VGND _0619_ _0658_ sg13g2_o21ai_1
X_5223_ _2132_ falu_i.falutop.data_in\[10\] _2133_ VPWR VGND sg13g2_xor2_1
X_5154_ falu_i.falutop.data_in\[11\] _2090_ _2091_ VPWR VGND sg13g2_nor2b_1
X_4105_ VGND VPWR net779 net952 _1108_ _1107_ sg13g2_a21oi_1
XFILLER_29_418 VPWR VGND sg13g2_decap_8
X_5085_ VPWR _2025_ _2024_ VGND sg13g2_inv_1
XFILLER_38_974 VPWR VGND sg13g2_decap_8
X_4036_ VGND VPWR _1059_ _1060_ _0222_ _1061_ sg13g2_a21oi_1
XFILLER_37_462 VPWR VGND sg13g2_decap_4
XFILLER_13_808 VPWR VGND sg13g2_decap_8
XFILLER_25_668 VPWR VGND sg13g2_decap_4
XFILLER_24_145 VPWR VGND sg13g2_fill_1
X_4938_ _1880_ _1881_ _1317_ _1882_ VPWR VGND sg13g2_nand3_1
X_4869_ _1814_ _1808_ _1812_ _1813_ VPWR VGND sg13g2_and3_1
XFILLER_21_896 VPWR VGND sg13g2_decap_8
XFILLER_21_67 VPWR VGND sg13g2_fill_2
XFILLER_43_1003 VPWR VGND sg13g2_decap_8
XFILLER_0_778 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_29_963 VPWR VGND sg13g2_decap_8
XFILLER_16_602 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_fill_2
XFILLER_44_944 VPWR VGND sg13g2_decap_8
XFILLER_24_690 VPWR VGND sg13g2_decap_8
XFILLER_31_649 VPWR VGND sg13g2_fill_1
XFILLER_12_874 VPWR VGND sg13g2_decap_8
XFILLER_8_867 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_35_977 VPWR VGND sg13g2_decap_8
XFILLER_21_115 VPWR VGND sg13g2_fill_1
X_2984_ ppwm_i.u_ppwm.u_mem.memory\[0\] _2310_ _2338_ VPWR VGND sg13g2_nor2_1
X_4723_ _1670_ _1246_ _1669_ VPWR VGND sg13g2_xnor2_1
X_4654_ _1602_ _1600_ _1601_ VPWR VGND sg13g2_nand2b_1
X_3605_ _0739_ net571 _0773_ _0774_ VPWR VGND sg13g2_a21o_1
X_4585_ _1534_ _1528_ _1532_ VPWR VGND sg13g2_xnor2_1
X_3536_ _2248_ net586 _0708_ VPWR VGND sg13g2_nor2_1
X_5206_ _2121_ falu_i.falutop.data_in\[4\] _2120_ VPWR VGND sg13g2_xnor2_1
X_3467_ _0643_ ppwm_i.u_ppwm.pwm_value\[0\] net608 VPWR VGND sg13g2_xnor2_1
X_3398_ VPWR VGND _2240_ _0575_ ppwm_i.u_ppwm.global_counter\[13\] _2239_ _0576_ ppwm_i.u_ppwm.global_counter\[14\]
+ sg13g2_a221oi_1
X_5137_ VGND VPWR _2071_ _2074_ _0309_ _2075_ sg13g2_a21oi_1
X_5068_ VGND VPWR _2007_ _2009_ _1983_ _1980_ sg13g2_a21oi_2
X_4019_ net805 VPWR _1047_ VGND falu_i.falutop.i2c_inst.state\[0\] _1046_ sg13g2_o21ai_1
XFILLER_26_944 VPWR VGND sg13g2_decap_8
XFILLER_16_56 VPWR VGND sg13g2_decap_4
XFILLER_13_627 VPWR VGND sg13g2_fill_2
XFILLER_41_969 VPWR VGND sg13g2_decap_8
XFILLER_32_11 VPWR VGND sg13g2_fill_2
X_5254__187 VPWR VGND net187 sg13g2_tiehi
XFILLER_21_682 VPWR VGND sg13g2_fill_2
XFILLER_32_55 VPWR VGND sg13g2_fill_1
XFILLER_10_1013 VPWR VGND sg13g2_decap_8
XFILLER_4_369 VPWR VGND sg13g2_fill_2
XFILLER_17_911 VPWR VGND sg13g2_decap_8
XFILLER_35_218 VPWR VGND sg13g2_fill_1
XFILLER_17_988 VPWR VGND sg13g2_decap_8
XFILLER_32_947 VPWR VGND sg13g2_decap_8
XFILLER_8_664 VPWR VGND sg13g2_fill_2
XFILLER_12_693 VPWR VGND sg13g2_decap_4
XFILLER_7_174 VPWR VGND sg13g2_fill_2
Xhold108 _1143_ VPWR VGND net480 sg13g2_dlygate4sd3_1
Xhold119 ppwm_i.u_ppwm.u_mem.memory\[63\] VPWR VGND net491 sg13g2_dlygate4sd3_1
X_4370_ VGND VPWR _1323_ _1321_ _1260_ sg13g2_or2_1
X_3321_ _0479_ _0500_ _0501_ VPWR VGND sg13g2_nor2_1
XFILLER_39_502 VPWR VGND sg13g2_decap_8
X_3252_ _0444_ net954 net1120 _0440_ VPWR VGND sg13g2_and3_1
X_3183_ _0397_ net512 ppwm_i.u_ppwm.u_mem.bit_count\[5\] VPWR VGND sg13g2_nand2_1
XFILLER_19_270 VPWR VGND sg13g2_fill_1
XFILLER_23_947 VPWR VGND sg13g2_decap_8
XFILLER_35_796 VPWR VGND sg13g2_fill_2
XFILLER_33_1002 VPWR VGND sg13g2_decap_8
XFILLER_34_295 VPWR VGND sg13g2_fill_1
X_2967_ net787 VPWR _2321_ VGND _2317_ _2320_ sg13g2_o21ai_1
X_5511__241 VPWR VGND net241 sg13g2_tiehi
X_2898_ VPWR _2252_ net376 VGND sg13g2_inv_1
X_4706_ _1653_ net738 net748 VPWR VGND sg13g2_nand2_2
X_4637_ _1404_ _1525_ net905 _1586_ VPWR VGND sg13g2_nand3_1
X_4568_ VPWR VGND _1373_ _1517_ _1508_ net631 _1518_ _1505_ sg13g2_a221oi_1
X_4499_ _1437_ _1438_ _1446_ _1449_ _1450_ VPWR VGND sg13g2_nor4_1
X_3519_ VGND VPWR _0688_ _0691_ _0692_ _0618_ sg13g2_a21oi_1
XFILLER_17_218 VPWR VGND sg13g2_fill_1
XFILLER_26_763 VPWR VGND sg13g2_fill_2
XFILLER_40_210 VPWR VGND sg13g2_fill_2
XFILLER_14_936 VPWR VGND sg13g2_decap_8
XFILLER_40_243 VPWR VGND sg13g2_fill_1
XFILLER_9_417 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_20_clk clknet_3_4__leaf_clk clknet_leaf_20_clk VPWR VGND sg13g2_buf_8
XFILLER_5_645 VPWR VGND sg13g2_fill_2
XFILLER_49_1020 VPWR VGND sg13g2_decap_8
XFILLER_4_15 VPWR VGND sg13g2_decap_8
XFILLER_4_188 VPWR VGND sg13g2_fill_1
XFILLER_4_26 VPWR VGND sg13g2_fill_1
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_49_866 VPWR VGND sg13g2_decap_8
XFILLER_1_1022 VPWR VGND sg13g2_decap_8
X_3870_ VGND VPWR _2197_ net645 _0154_ _0963_ sg13g2_a21oi_1
XFILLER_32_755 VPWR VGND sg13g2_fill_2
XFILLER_32_777 VPWR VGND sg13g2_decap_8
X_2821_ VPWR _2175_ net878 VGND sg13g2_inv_1
XFILLER_9_951 VPWR VGND sg13g2_decap_8
X_5540_ net60 VGND VPWR _0299_ falu_i.falutop.i2c_inst.result\[4\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_11_clk clknet_3_3__leaf_clk clknet_leaf_11_clk VPWR VGND sg13g2_buf_8
X_5471_ net343 VGND VPWR net973 falu_i.falutop.data_in\[2\] clknet_leaf_7_clk sg13g2_dfrbpq_2
X_4422_ _1374_ _2299_ _1303_ VPWR VGND sg13g2_nand2_2
X_4353_ _1304_ _1305_ _1306_ VPWR VGND sg13g2_nor2b_2
X_3304_ _0485_ net791 _2418_ VPWR VGND sg13g2_xnor2_1
X_4284_ _1237_ net729 net752 VPWR VGND sg13g2_nand2_2
X_3235_ _0433_ net1145 _0431_ VPWR VGND sg13g2_nand2_2
XFILLER_27_505 VPWR VGND sg13g2_fill_1
X_3166_ VGND VPWR _2287_ net681 _0025_ _0388_ sg13g2_a21oi_1
X_3097_ _2446_ _2433_ _2445_ VPWR VGND sg13g2_nand2_2
XFILLER_23_744 VPWR VGND sg13g2_decap_8
X_3999_ net1186 VPWR _1032_ VGND net883 _1021_ sg13g2_o21ai_1
Xhold472 falu_i.falutop.div_inst.rem\[4\] VPWR VGND net1124 sg13g2_dlygate4sd3_1
Xhold450 _0324_ VPWR VGND net1102 sg13g2_dlygate4sd3_1
Xhold461 _0034_ VPWR VGND net1113 sg13g2_dlygate4sd3_1
Xhold494 _0434_ VPWR VGND net1146 sg13g2_dlygate4sd3_1
Xhold483 falu_i.falutop.data_in\[3\] VPWR VGND net1135 sg13g2_dlygate4sd3_1
XFILLER_49_118 VPWR VGND sg13g2_fill_1
XFILLER_38_65 VPWR VGND sg13g2_fill_1
XFILLER_18_527 VPWR VGND sg13g2_decap_8
XFILLER_33_519 VPWR VGND sg13g2_decap_4
XFILLER_14_766 VPWR VGND sg13g2_decap_8
XFILLER_9_236 VPWR VGND sg13g2_fill_2
XFILLER_10_950 VPWR VGND sg13g2_decap_8
XFILLER_6_976 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_5_497 VPWR VGND sg13g2_fill_1
XFILLER_1_681 VPWR VGND sg13g2_fill_2
X_3020_ _2367_ net786 _2373_ _2374_ VPWR VGND sg13g2_a21o_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk clknet_leaf_0_clk VPWR VGND sg13g2_buf_8
X_5501__273 VPWR VGND net273 sg13g2_tiehi
X_4971_ _1914_ _1902_ _1912_ VPWR VGND sg13g2_xnor2_1
X_3922_ VGND VPWR _2177_ net677 _0180_ _0989_ sg13g2_a21oi_1
XFILLER_17_593 VPWR VGND sg13g2_fill_1
X_3853_ net826 VPWR _0955_ VGND net530 net658 sg13g2_o21ai_1
XFILLER_32_574 VPWR VGND sg13g2_fill_1
XFILLER_20_758 VPWR VGND sg13g2_decap_8
X_2804_ VPWR _2158_ net461 VGND sg13g2_inv_1
X_3784_ VGND VPWR _2226_ net655 _0111_ _0920_ sg13g2_a21oi_1
X_5523_ net182 VGND VPWR net436 falu_i.falutop.div_inst.quo\[3\] clknet_leaf_41_clk
+ sg13g2_dfrbpq_1
X_5454_ net70 VGND VPWR _0213_ ppwm_i.u_ppwm.u_mem.bit_count\[1\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_5385_ net282 VGND VPWR _0144_ ppwm_i.u_ppwm.u_mem.memory\[44\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4405_ _1355_ _1354_ _1357_ VPWR VGND sg13g2_xor2_1
X_4336_ net716 net710 _1286_ _1289_ VPWR VGND sg13g2_nor3_2
XFILLER_8_1028 VPWR VGND sg13g2_fill_1
X_5312__77 VPWR VGND net77 sg13g2_tiehi
X_4267_ _1220_ net745 net769 VPWR VGND sg13g2_nand2_2
X_3218_ ppwm_i.u_ppwm.u_pwm.counter\[8\] ppwm_i.u_ppwm.u_pwm.counter\[7\] ppwm_i.u_ppwm.u_pwm.counter\[9\]
+ _0422_ VPWR VGND ppwm_i.u_ppwm.u_pwm.counter\[6\] sg13g2_nand4_1
X_4198_ _1170_ net567 _1169_ VPWR VGND sg13g2_nand2_1
XFILLER_39_184 VPWR VGND sg13g2_decap_8
X_3149_ VGND VPWR net802 _0376_ _0019_ _0377_ sg13g2_a21oi_1
XFILLER_43_806 VPWR VGND sg13g2_fill_2
X_5536__96 VPWR VGND net96 sg13g2_tiehi
XFILLER_40_99 VPWR VGND sg13g2_fill_2
XFILLER_3_924 VPWR VGND sg13g2_decap_8
Xhold280 _0292_ VPWR VGND net932 sg13g2_dlygate4sd3_1
XFILLER_49_64 VPWR VGND sg13g2_decap_8
Xhold291 _0424_ VPWR VGND net943 sg13g2_dlygate4sd3_1
Xfanout760 falu_i.falutop.alu_data_in\[3\] net760 VPWR VGND sg13g2_buf_8
Xfanout782 ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] net782 VPWR VGND sg13g2_buf_8
Xfanout793 ppwm_i.u_ppwm.pc\[0\] net793 VPWR VGND sg13g2_buf_8
XFILLER_19_814 VPWR VGND sg13g2_decap_8
Xfanout771 net964 net771 VPWR VGND sg13g2_buf_8
XFILLER_46_666 VPWR VGND sg13g2_fill_2
XFILLER_45_132 VPWR VGND sg13g2_fill_2
XFILLER_14_552 VPWR VGND sg13g2_fill_2
X_5542__44 VPWR VGND net44 sg13g2_tiehi
XFILLER_46_4 VPWR VGND sg13g2_fill_1
X_5170_ VGND VPWR _2304_ net620 _0314_ _2103_ sg13g2_a21oi_1
X_4121_ _1122_ _1121_ _1114_ _1123_ VPWR VGND sg13g2_a21o_1
X_4052_ _2291_ falu_i.falutop.i2c_inst.op\[1\] _2292_ _2293_ _1073_ VPWR VGND sg13g2_nor4_1
XFILLER_49_482 VPWR VGND sg13g2_decap_8
X_3003_ _2357_ net689 ppwm_i.u_ppwm.u_mem.memory\[37\] net696 ppwm_i.u_ppwm.u_mem.memory\[30\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_633 VPWR VGND sg13g2_fill_1
XFILLER_37_622 VPWR VGND sg13g2_decap_8
Xinput4 ui_in[4] net4 VPWR VGND sg13g2_buf_1
XFILLER_40_809 VPWR VGND sg13g2_fill_2
X_4954_ _1897_ _1896_ _1895_ VPWR VGND sg13g2_nand2b_1
XFILLER_17_390 VPWR VGND sg13g2_fill_2
XFILLER_36_198 VPWR VGND sg13g2_decap_8
X_3905_ net834 VPWR _0981_ VGND net482 net669 sg13g2_o21ai_1
X_4885_ net615 VPWR _1830_ VGND _1788_ _1828_ sg13g2_o21ai_1
X_3836_ VGND VPWR _2209_ net643 _0137_ _0946_ sg13g2_a21oi_1
X_3767_ net827 VPWR _0912_ VGND ppwm_i.u_ppwm.u_mem.memory\[3\] net659 sg13g2_o21ai_1
X_5506_ net261 VGND VPWR net941 falu_i.falutop.div_inst.val\[1\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_2
X_3698_ VGND VPWR _0857_ _0858_ _0859_ _0618_ sg13g2_a21oi_1
XFILLER_10_14 VPWR VGND sg13g2_fill_1
X_5437_ net143 VGND VPWR net533 ppwm_i.u_ppwm.u_mem.memory\[96\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_5368_ net316 VGND VPWR net960 ppwm_i.u_ppwm.u_mem.memory\[27\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_5299_ net99 VGND VPWR _0061_ ppwm_i.u_ppwm.global_counter\[16\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
X_4319_ VGND VPWR _1270_ _1271_ _1272_ _1217_ sg13g2_a21oi_1
X_5404__244 VPWR VGND net244 sg13g2_tiehi
XFILLER_15_305 VPWR VGND sg13g2_fill_2
XFILLER_16_839 VPWR VGND sg13g2_decap_8
XFILLER_43_647 VPWR VGND sg13g2_fill_2
XFILLER_24_872 VPWR VGND sg13g2_decap_8
XFILLER_38_419 VPWR VGND sg13g2_fill_2
Xfanout590 _0610_ net590 VPWR VGND sg13g2_buf_8
XFILLER_18_8 VPWR VGND sg13g2_fill_1
XFILLER_19_633 VPWR VGND sg13g2_fill_2
XFILLER_47_953 VPWR VGND sg13g2_decap_8
XFILLER_33_124 VPWR VGND sg13g2_fill_2
XFILLER_15_861 VPWR VGND sg13g2_decap_8
X_4670_ VGND VPWR net631 _1610_ _1618_ _1617_ sg13g2_a21oi_1
X_3621_ _0678_ _0714_ _0789_ VPWR VGND sg13g2_nor2_1
X_3552_ VGND VPWR net974 net593 _0724_ _0723_ sg13g2_a21oi_1
X_3483_ _0658_ net785 net611 VPWR VGND sg13g2_xnor2_1
X_5222_ net776 VPWR _2132_ VGND falu_i.falutop.data_in\[8\] falu_i.falutop.data_in\[9\]
+ sg13g2_o21ai_1
X_5153_ falu_i.falutop.data_in\[8\] falu_i.falutop.data_in\[9\] falu_i.falutop.data_in\[10\]
+ _2090_ VPWR VGND sg13g2_nor3_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
X_4104_ net779 net396 _1107_ VPWR VGND sg13g2_nor2b_1
X_5084_ _1804_ VPWR _2024_ VGND _1652_ _1949_ sg13g2_o21ai_1
XFILLER_49_290 VPWR VGND sg13g2_decap_8
XFILLER_38_953 VPWR VGND sg13g2_decap_8
X_4035_ net804 VPWR _1061_ VGND net1043 _1059_ sg13g2_o21ai_1
XFILLER_36_1011 VPWR VGND sg13g2_decap_8
X_4937_ _1829_ _1879_ _1827_ _1881_ VPWR VGND sg13g2_nand3_1
X_4868_ _1752_ VPWR _1813_ VGND _1809_ _1811_ sg13g2_o21ai_1
XFILLER_21_875 VPWR VGND sg13g2_decap_8
X_3819_ net831 VPWR _0938_ VGND ppwm_i.u_ppwm.u_mem.memory\[30\] net643 sg13g2_o21ai_1
X_4799_ _1743_ _1744_ _1745_ VPWR VGND sg13g2_nor2_1
X_5287__123 VPWR VGND net123 sg13g2_tiehi
XFILLER_0_757 VPWR VGND sg13g2_decap_8
XFILLER_29_942 VPWR VGND sg13g2_decap_8
XFILLER_44_923 VPWR VGND sg13g2_decap_8
XFILLER_12_853 VPWR VGND sg13g2_decap_8
XFILLER_8_846 VPWR VGND sg13g2_decap_8
XFILLER_7_356 VPWR VGND sg13g2_decap_4
XFILLER_3_551 VPWR VGND sg13g2_fill_1
XFILLER_11_90 VPWR VGND sg13g2_fill_2
XFILLER_4_1020 VPWR VGND sg13g2_decap_8
XFILLER_19_463 VPWR VGND sg13g2_decap_8
XFILLER_35_956 VPWR VGND sg13g2_decap_8
X_2983_ VGND VPWR _2335_ _2336_ _2337_ _2254_ sg13g2_a21oi_1
X_4722_ _1215_ VPWR _1669_ VGND _1218_ _1611_ sg13g2_o21ai_1
X_4653_ VGND VPWR _1537_ _1538_ _1601_ _1540_ sg13g2_a21oi_1
X_3604_ _0649_ _0770_ _0771_ _0772_ _0773_ VPWR VGND sg13g2_nor4_1
X_4584_ _1533_ _1532_ _1528_ VPWR VGND sg13g2_nand2b_1
X_3535_ VPWR VGND _0707_ net798 _0693_ _2249_ _0075_ net572 sg13g2_a221oi_1
X_3466_ VGND VPWR net589 _0640_ _0642_ _0641_ sg13g2_a21oi_1
X_5205_ _2097_ net777 _2120_ VPWR VGND sg13g2_nor2b_1
X_3397_ VGND VPWR ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] _2264_ _0575_ _0574_ sg13g2_a21oi_1
X_5136_ net815 VPWR _2075_ VGND net1071 net627 sg13g2_o21ai_1
X_5067_ _1983_ _2007_ _1980_ _2008_ VPWR VGND sg13g2_nand3_1
X_4018_ net2 net1 _1046_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_923 VPWR VGND sg13g2_decap_8
XFILLER_37_271 VPWR VGND sg13g2_fill_2
XFILLER_41_948 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_fill_1
XFILLER_12_138 VPWR VGND sg13g2_decap_8
XFILLER_21_661 VPWR VGND sg13g2_fill_1
XFILLER_20_193 VPWR VGND sg13g2_fill_1
XFILLER_5_816 VPWR VGND sg13g2_decap_4
XFILLER_4_359 VPWR VGND sg13g2_decap_4
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_28_282 VPWR VGND sg13g2_decap_8
XFILLER_29_794 VPWR VGND sg13g2_fill_2
XFILLER_44_753 VPWR VGND sg13g2_fill_2
XFILLER_17_967 VPWR VGND sg13g2_decap_8
XFILLER_32_904 VPWR VGND sg13g2_fill_2
XFILLER_43_274 VPWR VGND sg13g2_fill_2
XFILLER_31_447 VPWR VGND sg13g2_fill_2
XFILLER_40_981 VPWR VGND sg13g2_decap_8
Xhold109 ppwm_i.u_ppwm.u_mem.memory\[36\] VPWR VGND net481 sg13g2_dlygate4sd3_1
XFILLER_7_197 VPWR VGND sg13g2_fill_2
X_3320_ net1162 _0495_ _0500_ VPWR VGND sg13g2_nor2_1
XFILLER_26_1021 VPWR VGND sg13g2_decap_8
X_3251_ VGND VPWR ppwm_i.u_ppwm.global_counter\[10\] _0440_ _0443_ net954 sg13g2_a21oi_1
X_3182_ VGND VPWR _2279_ net683 _0033_ _0396_ sg13g2_a21oi_1
XFILLER_34_241 VPWR VGND sg13g2_decap_8
XFILLER_23_926 VPWR VGND sg13g2_decap_8
XFILLER_34_274 VPWR VGND sg13g2_fill_2
X_2966_ _2320_ _2318_ _2319_ VPWR VGND sg13g2_nand2_1
X_4705_ _1652_ net711 net750 VPWR VGND sg13g2_nand2_1
XFILLER_30_480 VPWR VGND sg13g2_fill_1
X_2897_ _2251_ net1165 VPWR VGND sg13g2_inv_2
X_4636_ VGND VPWR _1404_ _1525_ _1585_ net905 sg13g2_a21oi_1
X_4567_ _1513_ _1514_ _1512_ _1517_ VPWR VGND _1516_ sg13g2_nand4_1
X_4498_ _1443_ _1445_ _1439_ _1449_ VPWR VGND _1448_ sg13g2_nand4_1
X_3518_ _0689_ _0690_ _0691_ VPWR VGND sg13g2_nor2b_1
X_3449_ _0625_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] net594 VPWR VGND sg13g2_nand2_1
X_5119_ _2026_ _2057_ _2058_ VPWR VGND sg13g2_nor2_1
XFILLER_14_915 VPWR VGND sg13g2_decap_8
XFILLER_26_753 VPWR VGND sg13g2_fill_1
XFILLER_43_55 VPWR VGND sg13g2_fill_1
XFILLER_22_992 VPWR VGND sg13g2_decap_8
XFILLER_49_801 VPWR VGND sg13g2_decap_8
XFILLER_48_311 VPWR VGND sg13g2_fill_2
XFILLER_48_300 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_49_845 VPWR VGND sg13g2_decap_8
XFILLER_0_384 VPWR VGND sg13g2_decap_8
XFILLER_0_395 VPWR VGND sg13g2_fill_1
XFILLER_1_1001 VPWR VGND sg13g2_decap_8
XFILLER_17_764 VPWR VGND sg13g2_fill_1
XFILLER_16_263 VPWR VGND sg13g2_fill_1
XFILLER_17_1009 VPWR VGND sg13g2_decap_8
XFILLER_31_222 VPWR VGND sg13g2_fill_1
XFILLER_9_930 VPWR VGND sg13g2_decap_8
X_2820_ VPWR _2174_ net510 VGND sg13g2_inv_1
XFILLER_12_491 VPWR VGND sg13g2_decap_4
XFILLER_13_992 VPWR VGND sg13g2_decap_8
X_5470_ net345 VGND VPWR net902 falu_i.falutop.data_in\[1\] clknet_leaf_8_clk sg13g2_dfrbpq_2
X_4421_ _2299_ _1303_ _1373_ VPWR VGND sg13g2_and2_1
X_5309__83 VPWR VGND net83 sg13g2_tiehi
X_4352_ net772 net771 _1305_ VPWR VGND sg13g2_nor2_1
X_5324__53 VPWR VGND net53 sg13g2_tiehi
X_5428__180 VPWR VGND net180 sg13g2_tiehi
X_3303_ VGND VPWR _2307_ _2310_ _0484_ net1162 sg13g2_a21oi_1
X_4283_ net729 net754 _1236_ VPWR VGND sg13g2_and2_1
X_3234_ _0431_ net1108 _0049_ VPWR VGND sg13g2_nor2_1
X_3165_ net807 VPWR _0388_ VGND net785 net681 sg13g2_o21ai_1
X_3096_ falu_i.falutop.i2c_inst.counter\[1\] falu_i.falutop.i2c_inst.counter\[0\]
+ _2445_ VPWR VGND sg13g2_nor2b_2
XFILLER_23_723 VPWR VGND sg13g2_decap_8
X_5435__151 VPWR VGND net151 sg13g2_tiehi
XFILLER_10_406 VPWR VGND sg13g2_fill_2
X_3998_ net1052 _1030_ _1031_ _0214_ VPWR VGND sg13g2_nor3_1
X_2949_ VPWR _2303_ net754 VGND sg13g2_inv_1
X_4619_ VGND VPWR _1496_ _1565_ _1568_ _1318_ sg13g2_a21oi_1
Xhold440 ppwm_i.u_ppwm.global_counter\[7\] VPWR VGND net1092 sg13g2_dlygate4sd3_1
Xhold451 falu_i.falutop.data_in\[12\] VPWR VGND net1103 sg13g2_dlygate4sd3_1
Xhold462 falu_i.falutop.data_in\[4\] VPWR VGND net1114 sg13g2_dlygate4sd3_1
Xhold473 ppwm_i.u_ppwm.global_counter\[16\] VPWR VGND net1125 sg13g2_dlygate4sd3_1
Xhold495 _0050_ VPWR VGND net1147 sg13g2_dlygate4sd3_1
Xhold484 _0316_ VPWR VGND net1136 sg13g2_dlygate4sd3_1
X_5442__122 VPWR VGND net122 sg13g2_tiehi
XFILLER_38_11 VPWR VGND sg13g2_fill_2
XFILLER_18_506 VPWR VGND sg13g2_fill_2
XFILLER_45_358 VPWR VGND sg13g2_fill_1
XFILLER_13_200 VPWR VGND sg13g2_decap_8
X_5414__224 VPWR VGND net224 sg13g2_tiehi
XFILLER_14_789 VPWR VGND sg13g2_fill_1
XFILLER_6_955 VPWR VGND sg13g2_decap_8
XFILLER_49_675 VPWR VGND sg13g2_decap_4
XFILLER_23_1024 VPWR VGND sg13g2_decap_4
XFILLER_49_697 VPWR VGND sg13g2_decap_8
XFILLER_36_303 VPWR VGND sg13g2_fill_2
XFILLER_24_509 VPWR VGND sg13g2_fill_1
X_4970_ _1913_ _1902_ _1912_ VPWR VGND sg13g2_nand2_1
X_3921_ net840 VPWR _0989_ VGND net886 net677 sg13g2_o21ai_1
X_3852_ VGND VPWR _2203_ net657 _0145_ _0954_ sg13g2_a21oi_1
XFILLER_20_726 VPWR VGND sg13g2_fill_1
X_2803_ VPWR _2157_ net559 VGND sg13g2_inv_1
X_5522_ net186 VGND VPWR net412 falu_i.falutop.div_inst.quo\[2\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_3783_ net824 VPWR _0920_ VGND net888 net655 sg13g2_o21ai_1
XFILLER_9_793 VPWR VGND sg13g2_fill_2
XFILLER_30_1028 VPWR VGND sg13g2_fill_1
X_5453_ net74 VGND VPWR net379 ppwm_i.u_ppwm.u_mem.bit_count\[0\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
X_5384_ net284 VGND VPWR _0143_ ppwm_i.u_ppwm.u_mem.memory\[43\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_4404_ _1356_ _1354_ _1355_ VPWR VGND sg13g2_nand2b_1
X_4335_ _1287_ _1284_ _1288_ VPWR VGND sg13g2_nor2b_2
XFILLER_8_1007 VPWR VGND sg13g2_decap_8
X_4266_ net744 net770 _1219_ VPWR VGND sg13g2_and2_1
X_4197_ _1169_ _1123_ _1124_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_815 VPWR VGND sg13g2_fill_1
X_3217_ ppwm_i.u_ppwm.u_pwm.counter\[0\] net809 ppwm_i.u_ppwm.u_pwm.counter\[1\] _0421_
+ VPWR VGND sg13g2_nand3_1
X_3148_ net804 VPWR _0377_ VGND net908 _0376_ sg13g2_o21ai_1
XFILLER_42_306 VPWR VGND sg13g2_decap_8
X_3079_ net985 net1013 _2430_ VPWR VGND sg13g2_nor2_2
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_236 VPWR VGND sg13g2_decap_8
XFILLER_11_759 VPWR VGND sg13g2_fill_1
XFILLER_3_903 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
Xhold270 ppwm_i.u_ppwm.u_mem.memory\[74\] VPWR VGND net922 sg13g2_dlygate4sd3_1
XFILLER_6_4 VPWR VGND sg13g2_fill_2
XFILLER_2_435 VPWR VGND sg13g2_fill_2
Xhold292 _0046_ VPWR VGND net944 sg13g2_dlygate4sd3_1
Xhold281 ppwm_i.u_ppwm.u_mem.memory\[13\] VPWR VGND net933 sg13g2_dlygate4sd3_1
Xfanout750 falu_i.falutop.alu_data_in\[5\] net750 VPWR VGND sg13g2_buf_8
Xfanout783 net1194 net783 VPWR VGND sg13g2_buf_1
Xfanout794 ppwm_i.u_ppwm.pc\[0\] net794 VPWR VGND sg13g2_buf_8
Xfanout761 net764 net761 VPWR VGND sg13g2_buf_2
Xfanout772 net938 net772 VPWR VGND sg13g2_buf_8
XFILLER_46_623 VPWR VGND sg13g2_fill_2
XFILLER_45_100 VPWR VGND sg13g2_fill_1
X_5297__103 VPWR VGND net103 sg13g2_tiehi
XFILLER_45_188 VPWR VGND sg13g2_fill_1
XFILLER_14_520 VPWR VGND sg13g2_fill_2
XFILLER_41_383 VPWR VGND sg13g2_decap_8
XFILLER_14_597 VPWR VGND sg13g2_decap_8
XFILLER_6_730 VPWR VGND sg13g2_fill_2
XFILLER_6_796 VPWR VGND sg13g2_decap_8
XFILLER_5_295 VPWR VGND sg13g2_fill_2
X_4120_ _1122_ falu_i.falutop.div_inst.b1\[3\] falu_i.falutop.div_inst.acc\[3\] VPWR
+ VGND sg13g2_xnor2_1
X_4051_ net797 _1072_ _0226_ VPWR VGND sg13g2_nor2_1
X_3002_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[2\] _2354_ net699 ppwm_i.u_ppwm.u_mem.memory\[23\]
+ _2356_ net701 sg13g2_a221oi_1
Xinput5 ui_in[5] net5 VPWR VGND sg13g2_buf_1
X_4953_ net733 net705 _1896_ VPWR VGND sg13g2_nor2_1
X_3904_ VGND VPWR _2185_ net647 _0171_ _0980_ sg13g2_a21oi_1
X_4884_ _1829_ _1788_ _1828_ VPWR VGND sg13g2_nand2_1
X_3835_ net829 VPWR _0946_ VGND ppwm_i.u_ppwm.u_mem.memory\[38\] net643 sg13g2_o21ai_1
XFILLER_20_556 VPWR VGND sg13g2_fill_2
X_3766_ VGND VPWR _2233_ net661 _0102_ _0911_ sg13g2_a21oi_1
XFILLER_9_590 VPWR VGND sg13g2_fill_1
X_5505_ net265 VGND VPWR _0264_ falu_i.falutop.div_inst.val\[0\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_2
X_5436_ net147 VGND VPWR _0195_ ppwm_i.u_ppwm.u_mem.memory\[95\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
X_3697_ VGND VPWR ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] net600 _0858_ _0850_ sg13g2_a21oi_1
XFILLER_0_939 VPWR VGND sg13g2_decap_8
X_5367_ net318 VGND VPWR _0126_ ppwm_i.u_ppwm.u_mem.memory\[26\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_5298_ net101 VGND VPWR _0060_ ppwm_i.u_ppwm.global_counter\[15\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
X_4318_ _1271_ net752 net729 VPWR VGND sg13g2_nand2b_1
X_4249_ _1208_ net494 _1105_ VPWR VGND sg13g2_nand2_1
XFILLER_19_35 VPWR VGND sg13g2_fill_1
XFILLER_42_136 VPWR VGND sg13g2_fill_1
XFILLER_15_339 VPWR VGND sg13g2_decap_8
XFILLER_24_851 VPWR VGND sg13g2_decap_8
XFILLER_11_545 VPWR VGND sg13g2_decap_8
XFILLER_3_733 VPWR VGND sg13g2_decap_4
X_5264__168 VPWR VGND net168 sg13g2_tiehi
XFILLER_47_932 VPWR VGND sg13g2_decap_8
Xfanout591 net592 net591 VPWR VGND sg13g2_buf_8
Xfanout580 _0608_ net580 VPWR VGND sg13g2_buf_8
XFILLER_46_486 VPWR VGND sg13g2_decap_8
XFILLER_46_453 VPWR VGND sg13g2_decap_4
XFILLER_19_689 VPWR VGND sg13g2_decap_8
XFILLER_34_615 VPWR VGND sg13g2_fill_2
XFILLER_46_497 VPWR VGND sg13g2_fill_1
XFILLER_15_840 VPWR VGND sg13g2_decap_8
XFILLER_33_147 VPWR VGND sg13g2_fill_1
XFILLER_42_692 VPWR VGND sg13g2_decap_8
X_3620_ _0624_ _0694_ _0788_ VPWR VGND sg13g2_nor2_1
X_3551_ _2270_ net593 _0723_ VPWR VGND sg13g2_nor2_1
X_3482_ _0657_ net785 net611 VPWR VGND sg13g2_nand2_1
XFILLER_44_2 VPWR VGND sg13g2_fill_1
X_5221_ net475 net625 _2131_ VPWR VGND sg13g2_nor2_1
X_5152_ VGND VPWR _2085_ _2088_ _0310_ _2089_ sg13g2_a21oi_1
X_4103_ _1106_ _1098_ _1104_ VPWR VGND sg13g2_nand2_2
X_5083_ _2023_ _2021_ _2022_ VPWR VGND sg13g2_nand2_2
X_4034_ _1050_ _1056_ _1060_ VPWR VGND sg13g2_nor2_1
XFILLER_40_607 VPWR VGND sg13g2_fill_2
XFILLER_24_136 VPWR VGND sg13g2_decap_8
XFILLER_40_629 VPWR VGND sg13g2_fill_2
X_4936_ _1829_ _1827_ _1879_ _1880_ VPWR VGND sg13g2_a21o_1
X_4867_ _1751_ _1810_ _1812_ VPWR VGND _1811_ sg13g2_nand3b_1
XFILLER_20_331 VPWR VGND sg13g2_decap_4
XFILLER_21_854 VPWR VGND sg13g2_decap_8
X_3818_ VGND VPWR _2214_ net660 _0128_ _0937_ sg13g2_a21oi_1
XFILLER_20_364 VPWR VGND sg13g2_decap_8
X_4798_ _1744_ net751 net738 net748 net742 VPWR VGND sg13g2_a22oi_1
XFILLER_21_69 VPWR VGND sg13g2_fill_1
X_3749_ net912 falu_i.falutop.i2c_inst.op\[1\] net686 _0093_ VPWR VGND sg13g2_mux2_1
X_5419_ net214 VGND VPWR net546 ppwm_i.u_ppwm.u_mem.memory\[78\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_28_431 VPWR VGND sg13g2_fill_2
XFILLER_29_998 VPWR VGND sg13g2_decap_8
XFILLER_16_637 VPWR VGND sg13g2_decap_8
XFILLER_44_979 VPWR VGND sg13g2_decap_8
XFILLER_15_147 VPWR VGND sg13g2_decap_4
XFILLER_31_618 VPWR VGND sg13g2_decap_8
XFILLER_12_810 VPWR VGND sg13g2_fill_2
XFILLER_12_832 VPWR VGND sg13g2_decap_8
XFILLER_3_585 VPWR VGND sg13g2_fill_2
XFILLER_30_8 VPWR VGND sg13g2_decap_4
XFILLER_38_206 VPWR VGND sg13g2_fill_1
X_2982_ VPWR VGND _2191_ net789 net691 _2196_ _2336_ net698 sg13g2_a221oi_1
X_4721_ _1668_ _1247_ _1273_ VPWR VGND sg13g2_xnor2_1
X_4652_ _1599_ _1591_ _1600_ VPWR VGND sg13g2_xor2_1
XFILLER_30_662 VPWR VGND sg13g2_fill_1
X_3603_ _0648_ _0714_ _0772_ VPWR VGND sg13g2_nor2_1
X_4583_ _1530_ _1531_ _1532_ VPWR VGND sg13g2_and2_1
X_3534_ _0702_ _0706_ _0707_ VPWR VGND sg13g2_and2_1
X_3465_ net579 VPWR _0641_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] net589 sg13g2_o21ai_1
X_5204_ net999 net623 _2119_ VPWR VGND sg13g2_nor2_1
X_3396_ _0574_ _0572_ _0573_ ppwm_i.u_ppwm.global_counter\[12\] _2241_ VPWR VGND sg13g2_a22oi_1
X_5135_ VGND VPWR net638 _2073_ _2074_ net630 sg13g2_a21oi_1
X_5066_ VPWR _2007_ _2006_ VGND sg13g2_inv_1
XFILLER_26_902 VPWR VGND sg13g2_decap_8
X_4017_ net796 _1044_ net935 _0219_ VPWR VGND sg13g2_nor3_1
XFILLER_16_25 VPWR VGND sg13g2_fill_1
XFILLER_16_36 VPWR VGND sg13g2_fill_1
XFILLER_16_69 VPWR VGND sg13g2_fill_1
XFILLER_25_445 VPWR VGND sg13g2_fill_2
XFILLER_26_979 VPWR VGND sg13g2_decap_8
XFILLER_41_927 VPWR VGND sg13g2_decap_8
XFILLER_34_990 VPWR VGND sg13g2_decap_8
XFILLER_40_437 VPWR VGND sg13g2_fill_1
X_4919_ _1860_ _1861_ _1857_ _1863_ VPWR VGND sg13g2_nand3_1
XFILLER_32_13 VPWR VGND sg13g2_fill_1
XFILLER_5_839 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_48_526 VPWR VGND sg13g2_fill_2
XFILLER_0_588 VPWR VGND sg13g2_decap_4
XFILLER_48_559 VPWR VGND sg13g2_fill_2
XFILLER_17_946 VPWR VGND sg13g2_decap_8
XFILLER_40_960 VPWR VGND sg13g2_decap_8
XFILLER_4_894 VPWR VGND sg13g2_decap_8
XFILLER_26_1000 VPWR VGND sg13g2_decap_8
X_3250_ net795 net1121 _0055_ VPWR VGND sg13g2_nor2_1
X_3181_ net810 VPWR _0396_ VGND ppwm_i.u_ppwm.pwm_value\[9\] net682 sg13g2_o21ai_1
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_23_905 VPWR VGND sg13g2_decap_8
X_2965_ _2319_ net695 _2185_ net703 _2180_ VPWR VGND sg13g2_a22oi_1
X_4704_ _1651_ net731 net715 VPWR VGND sg13g2_nand2_1
XFILLER_31_982 VPWR VGND sg13g2_decap_8
X_2896_ _2250_ ppwm_i.u_ppwm.pwm_value\[2\] VPWR VGND sg13g2_inv_2
X_4635_ net819 VPWR _1584_ VGND net1083 net628 sg13g2_o21ai_1
XFILLER_8_81 VPWR VGND sg13g2_decap_8
X_4566_ net640 _1515_ _1516_ VPWR VGND sg13g2_nor2_1
X_3517_ _0690_ _2249_ net586 VPWR VGND sg13g2_nand2_1
X_4497_ VPWR VGND _1226_ _1447_ _1324_ _1230_ _1448_ _1322_ sg13g2_a221oi_1
X_3448_ _0623_ VPWR _0624_ VGND _2248_ net594 sg13g2_o21ai_1
X_3379_ _0556_ VPWR _0557_ VGND _2241_ ppwm_i.u_ppwm.global_counter\[2\] sg13g2_o21ai_1
X_5118_ _2057_ _2024_ _2056_ VPWR VGND sg13g2_xnor2_1
X_5049_ _1988_ _1989_ _1990_ VPWR VGND sg13g2_nor2_1
XFILLER_25_242 VPWR VGND sg13g2_decap_4
XFILLER_26_776 VPWR VGND sg13g2_fill_2
XFILLER_41_757 VPWR VGND sg13g2_fill_2
XFILLER_40_234 VPWR VGND sg13g2_decap_8
XFILLER_13_426 VPWR VGND sg13g2_fill_2
XFILLER_13_448 VPWR VGND sg13g2_decap_4
XFILLER_22_971 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_49_824 VPWR VGND sg13g2_fill_2
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_36_529 VPWR VGND sg13g2_fill_2
XFILLER_16_231 VPWR VGND sg13g2_decap_4
XFILLER_31_234 VPWR VGND sg13g2_decap_8
XFILLER_13_971 VPWR VGND sg13g2_decap_8
XFILLER_12_481 VPWR VGND sg13g2_fill_2
XFILLER_31_289 VPWR VGND sg13g2_fill_1
XFILLER_9_986 VPWR VGND sg13g2_decap_8
X_4420_ _1372_ _1288_ _1338_ _1371_ VPWR VGND sg13g2_and3_1
X_4351_ _1304_ falu_i.falutop.alu_inst.op\[0\] VPWR VGND falu_i.falutop.alu_inst.op\[1\]
+ sg13g2_nand2b_2
X_3302_ VPWR VGND _0483_ net799 net1163 _2255_ _0066_ _2257_ sg13g2_a221oi_1
X_4282_ _1235_ _1233_ VPWR VGND _1231_ sg13g2_nand2b_2
XFILLER_39_301 VPWR VGND sg13g2_fill_2
X_3233_ net812 VPWR _0432_ VGND net1107 _0430_ sg13g2_o21ai_1
XFILLER_39_323 VPWR VGND sg13g2_decap_4
X_3164_ VGND VPWR _2288_ net681 _0024_ _0387_ sg13g2_a21oi_1
XFILLER_39_378 VPWR VGND sg13g2_fill_2
X_3095_ VGND VPWR net802 _2443_ _0004_ _2444_ sg13g2_a21oi_1
XFILLER_23_713 VPWR VGND sg13g2_fill_1
XFILLER_22_234 VPWR VGND sg13g2_fill_1
XFILLER_22_245 VPWR VGND sg13g2_fill_1
XFILLER_23_779 VPWR VGND sg13g2_decap_8
X_3997_ net808 VPWR _1031_ VGND net1051 _1025_ sg13g2_o21ai_1
X_2948_ VPWR _2302_ falu_i.falutop.alu_data_in\[7\] VGND sg13g2_inv_1
X_4618_ _1567_ _1496_ _1565_ VPWR VGND sg13g2_nand2_1
X_2879_ VPWR _2233_ net852 VGND sg13g2_inv_1
Xhold441 _0437_ VPWR VGND net1093 sg13g2_dlygate4sd3_1
XFILLER_2_628 VPWR VGND sg13g2_decap_8
Xhold452 _0325_ VPWR VGND net1104 sg13g2_dlygate4sd3_1
Xhold463 _0317_ VPWR VGND net1115 sg13g2_dlygate4sd3_1
X_4549_ VPWR VGND _1288_ _1289_ _1366_ net716 _1499_ _1294_ sg13g2_a221oi_1
Xhold430 _0329_ VPWR VGND net1082 sg13g2_dlygate4sd3_1
Xhold474 _0453_ VPWR VGND net1126 sg13g2_dlygate4sd3_1
Xhold485 falu_i.falutop.data_in\[7\] VPWR VGND net1137 sg13g2_dlygate4sd3_1
Xhold496 falu_i.falutop.data_in\[0\] VPWR VGND net1148 sg13g2_dlygate4sd3_1
XFILLER_26_595 VPWR VGND sg13g2_decap_8
XFILLER_9_205 VPWR VGND sg13g2_decap_8
XFILLER_9_238 VPWR VGND sg13g2_fill_1
XFILLER_16_1021 VPWR VGND sg13g2_decap_8
XFILLER_6_934 VPWR VGND sg13g2_decap_8
XFILLER_10_985 VPWR VGND sg13g2_decap_8
XFILLER_5_477 VPWR VGND sg13g2_decap_4
XFILLER_23_1003 VPWR VGND sg13g2_decap_8
XFILLER_37_838 VPWR VGND sg13g2_fill_1
XFILLER_36_326 VPWR VGND sg13g2_decap_8
X_3920_ VGND VPWR _2179_ net647 _0179_ _0988_ sg13g2_a21oi_1
XFILLER_44_381 VPWR VGND sg13g2_fill_2
X_5274__148 VPWR VGND net148 sg13g2_tiehi
X_3851_ net829 VPWR _0954_ VGND ppwm_i.u_ppwm.u_mem.memory\[45\] net657 sg13g2_o21ai_1
X_2802_ VPWR _2156_ net951 VGND sg13g2_inv_1
X_3782_ VGND VPWR _2227_ net660 _0110_ _0919_ sg13g2_a21oi_1
X_5521_ net190 VGND VPWR net400 falu_i.falutop.div_inst.quo\[1\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
XFILLER_30_1007 VPWR VGND sg13g2_decap_8
X_5452_ net78 VGND VPWR _0211_ ppwm_i.u_ppwm.u_mem.memory\[111\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_5383_ net286 VGND VPWR net855 ppwm_i.u_ppwm.u_mem.memory\[42\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4403_ VGND VPWR _1222_ _1255_ _1355_ _1254_ sg13g2_a21oi_1
X_4334_ _1285_ _1286_ _1287_ VPWR VGND sg13g2_nor2_1
X_4265_ VGND VPWR _1218_ _1216_ _1214_ sg13g2_or2_1
X_3216_ VGND VPWR _2273_ _0418_ _0043_ _0420_ sg13g2_a21oi_1
X_4196_ VGND VPWR net633 _1167_ _0275_ _1168_ sg13g2_a21oi_1
X_3147_ _2434_ net1007 _0376_ VPWR VGND sg13g2_nor2_1
XFILLER_43_808 VPWR VGND sg13g2_fill_1
XFILLER_27_337 VPWR VGND sg13g2_fill_2
X_3078_ _2427_ VPWR _0002_ VGND _2428_ _2429_ sg13g2_o21ai_1
XFILLER_46_1014 VPWR VGND sg13g2_decap_8
Xhold271 _0173_ VPWR VGND net923 sg13g2_dlygate4sd3_1
XFILLER_3_959 VPWR VGND sg13g2_decap_8
Xhold260 falu_i.falutop.i2c_inst.data_in\[17\] VPWR VGND net912 sg13g2_dlygate4sd3_1
XFILLER_2_469 VPWR VGND sg13g2_fill_2
Xhold293 falu_i.falutop.i2c_inst.data_in\[10\] VPWR VGND net945 sg13g2_dlygate4sd3_1
Xhold282 ppwm_i.u_ppwm.u_mem.data_sync2 VPWR VGND net934 sg13g2_dlygate4sd3_1
Xfanout751 falu_i.falutop.alu_data_in\[5\] net751 VPWR VGND sg13g2_buf_8
Xfanout740 falu_i.falutop.alu_data_in\[9\] net740 VPWR VGND sg13g2_buf_8
Xfanout773 net774 net773 VPWR VGND sg13g2_buf_2
Xfanout762 net763 net762 VPWR VGND sg13g2_buf_2
Xfanout784 net785 net784 VPWR VGND sg13g2_buf_8
XFILLER_46_602 VPWR VGND sg13g2_decap_8
XFILLER_19_849 VPWR VGND sg13g2_decap_8
Xfanout795 net796 net795 VPWR VGND sg13g2_buf_8
XFILLER_45_112 VPWR VGND sg13g2_decap_8
XFILLER_27_860 VPWR VGND sg13g2_fill_2
XFILLER_14_587 VPWR VGND sg13g2_decap_4
XFILLER_6_764 VPWR VGND sg13g2_fill_2
XFILLER_5_263 VPWR VGND sg13g2_decap_8
X_5529__153 VPWR VGND net153 sg13g2_tiehi
XFILLER_2_981 VPWR VGND sg13g2_decap_8
X_4050_ _1072_ _1071_ net1016 _1057_ _1046_ VPWR VGND sg13g2_a22oi_1
XFILLER_49_462 VPWR VGND sg13g2_decap_8
X_5302__90 VPWR VGND net90 sg13g2_tiehi
X_3001_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[9\] net689 _2355_ net789 sg13g2_a21oi_1
X_4952_ _1895_ net727 net748 VPWR VGND sg13g2_nand2_1
XFILLER_18_893 VPWR VGND sg13g2_decap_8
X_3903_ net834 VPWR _0980_ VGND net482 net646 sg13g2_o21ai_1
X_4883_ _1826_ _1789_ _1828_ VPWR VGND sg13g2_xor2_1
XFILLER_17_392 VPWR VGND sg13g2_fill_1
XFILLER_32_340 VPWR VGND sg13g2_decap_8
XFILLER_33_874 VPWR VGND sg13g2_decap_8
X_3834_ VGND VPWR _2209_ net664 _0136_ _0945_ sg13g2_a21oi_1
XFILLER_20_502 VPWR VGND sg13g2_fill_2
X_3765_ net828 VPWR _0911_ VGND ppwm_i.u_ppwm.u_mem.memory\[2\] net661 sg13g2_o21ai_1
X_3696_ VPWR _0857_ _0856_ VGND sg13g2_inv_1
X_5504_ net267 VGND VPWR _0263_ falu_i.falutop.div_inst.busy clknet_leaf_44_clk sg13g2_dfrbpq_1
X_5435_ net151 VGND VPWR _0194_ ppwm_i.u_ppwm.u_mem.memory\[94\] clknet_leaf_28_clk
+ sg13g2_dfrbpq_1
XFILLER_0_918 VPWR VGND sg13g2_decap_8
X_5366_ net320 VGND VPWR net509 ppwm_i.u_ppwm.u_mem.memory\[25\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_5297_ net103 VGND VPWR net976 ppwm_i.u_ppwm.global_counter\[14\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
X_4317_ _1269_ _1263_ _1239_ _1270_ VPWR VGND sg13g2_a21o_1
X_4248_ _1207_ VPWR _0288_ VGND _1098_ _1159_ sg13g2_o21ai_1
XFILLER_19_58 VPWR VGND sg13g2_decap_4
X_4179_ _1154_ net1009 _1155_ VPWR VGND sg13g2_xor2_1
XFILLER_15_307 VPWR VGND sg13g2_fill_1
XFILLER_24_830 VPWR VGND sg13g2_decap_8
XFILLER_23_351 VPWR VGND sg13g2_decap_8
Xclkbuf_3_3__f_clk clknet_0_clk clknet_3_3__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_11_579 VPWR VGND sg13g2_decap_8
XFILLER_13_1013 VPWR VGND sg13g2_decap_8
XFILLER_3_712 VPWR VGND sg13g2_decap_8
XFILLER_3_789 VPWR VGND sg13g2_decap_8
XFILLER_3_756 VPWR VGND sg13g2_decap_4
XFILLER_2_244 VPWR VGND sg13g2_decap_4
XFILLER_2_266 VPWR VGND sg13g2_fill_1
XFILLER_47_911 VPWR VGND sg13g2_decap_8
Xfanout581 net583 net581 VPWR VGND sg13g2_buf_8
Xfanout570 _0814_ net570 VPWR VGND sg13g2_buf_8
Xfanout592 net593 net592 VPWR VGND sg13g2_buf_8
X_5559__157 VPWR VGND net157 sg13g2_tiehi
XFILLER_19_657 VPWR VGND sg13g2_decap_4
XFILLER_20_1028 VPWR VGND sg13g2_fill_1
XFILLER_47_988 VPWR VGND sg13g2_decap_8
XFILLER_15_896 VPWR VGND sg13g2_decap_8
XFILLER_30_866 VPWR VGND sg13g2_decap_4
X_3550_ _0721_ VPWR _0722_ VGND _0715_ _0717_ sg13g2_o21ai_1
X_5220_ _2128_ VPWR _0337_ VGND net622 _2130_ sg13g2_o21ai_1
X_3481_ VPWR VGND net571 _0652_ _0655_ _0622_ _0656_ _0648_ sg13g2_a221oi_1
X_5151_ net815 VPWR _2089_ VGND net1029 net627 sg13g2_o21ai_1
X_5243__209 VPWR VGND net209 sg13g2_tiehi
X_5082_ _1944_ _1947_ _1987_ _2022_ VPWR VGND sg13g2_or3_1
X_4102_ _1097_ _1103_ _1105_ VPWR VGND sg13g2_nor2_2
XFILLER_38_933 VPWR VGND sg13g2_fill_2
XFILLER_38_922 VPWR VGND sg13g2_decap_8
X_4033_ _1059_ _1058_ VPWR VGND _1057_ sg13g2_nand2b_2
XFILLER_38_988 VPWR VGND sg13g2_decap_8
XFILLER_25_616 VPWR VGND sg13g2_fill_2
XFILLER_37_498 VPWR VGND sg13g2_decap_4
X_4935_ _1876_ _1841_ _1879_ VPWR VGND sg13g2_xor2_1
X_4866_ _1811_ net755 net723 net761 net718 VPWR VGND sg13g2_a22oi_1
XFILLER_21_833 VPWR VGND sg13g2_decap_8
X_3817_ net829 VPWR _0937_ VGND net959 net660 sg13g2_o21ai_1
X_4797_ _1653_ _1687_ _1743_ VPWR VGND sg13g2_nor2_1
X_3748_ VGND VPWR _2291_ net685 _0092_ _0903_ sg13g2_a21oi_1
XFILLER_4_509 VPWR VGND sg13g2_decap_4
X_3679_ _0842_ _0838_ _0841_ VPWR VGND sg13g2_xnor2_1
X_5418_ net216 VGND VPWR net552 ppwm_i.u_ppwm.u_mem.memory\[77\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_5349_ net354 VGND VPWR net442 ppwm_i.u_ppwm.u_mem.memory\[8\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_43_1028 VPWR VGND sg13g2_fill_1
XFILLER_43_1017 VPWR VGND sg13g2_decap_8
XFILLER_29_977 VPWR VGND sg13g2_decap_8
XFILLER_44_958 VPWR VGND sg13g2_decap_8
XFILLER_16_649 VPWR VGND sg13g2_decap_8
XFILLER_43_457 VPWR VGND sg13g2_fill_1
XFILLER_24_671 VPWR VGND sg13g2_decap_8
XFILLER_7_303 VPWR VGND sg13g2_decap_8
XFILLER_12_888 VPWR VGND sg13g2_decap_8
XFILLER_7_336 VPWR VGND sg13g2_decap_8
X_5385__282 VPWR VGND net282 sg13g2_tiehi
XFILLER_39_708 VPWR VGND sg13g2_decap_4
XFILLER_23_8 VPWR VGND sg13g2_decap_8
XFILLER_47_796 VPWR VGND sg13g2_fill_2
XFILLER_34_402 VPWR VGND sg13g2_decap_8
X_2981_ _2335_ net695 _2186_ net703 _2181_ VPWR VGND sg13g2_a22oi_1
XFILLER_15_660 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_41_clk clknet_3_1__leaf_clk clknet_leaf_41_clk VPWR VGND sg13g2_buf_8
X_4720_ _1246_ _1273_ _1667_ VPWR VGND sg13g2_nor2_1
X_4651_ _1597_ _1536_ _1599_ VPWR VGND sg13g2_xor2_1
XFILLER_30_652 VPWR VGND sg13g2_fill_1
X_3602_ _0626_ _0694_ _0771_ VPWR VGND sg13g2_nor2_1
X_4582_ net717 net736 net754 _1531_ VPWR VGND sg13g2_a21o_1
XFILLER_7_881 VPWR VGND sg13g2_decap_8
X_3533_ VGND VPWR net577 _0705_ _0706_ net572 sg13g2_a21oi_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
X_3464_ VGND VPWR ppwm_i.u_ppwm.global_counter\[10\] net595 _0640_ _0639_ sg13g2_a21oi_1
X_5203_ VGND VPWR net623 _2118_ _0332_ _2116_ sg13g2_a21oi_1
X_5134_ _2073_ falu_i.falutop.div_inst.rem\[6\] _2072_ VPWR VGND sg13g2_xnor2_1
X_3395_ _0573_ _2266_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] _2265_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\]
+ VPWR VGND sg13g2_a22oi_1
X_5065_ _2006_ _1984_ _2004_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_229 VPWR VGND sg13g2_decap_8
XFILLER_38_752 VPWR VGND sg13g2_decap_8
X_4016_ VGND VPWR net934 _0906_ _1045_ net883 sg13g2_a21oi_1
XFILLER_26_958 VPWR VGND sg13g2_decap_8
XFILLER_40_416 VPWR VGND sg13g2_decap_8
XFILLER_12_107 VPWR VGND sg13g2_decap_8
X_4918_ _1862_ _1857_ _1860_ _1861_ VPWR VGND sg13g2_and3_1
Xclkbuf_leaf_32_clk clknet_3_7__leaf_clk clknet_leaf_32_clk VPWR VGND sg13g2_buf_8
XFILLER_33_490 VPWR VGND sg13g2_decap_8
X_4849_ net742 net706 _1653_ _1794_ VPWR VGND sg13g2_nor3_1
XFILLER_4_306 VPWR VGND sg13g2_fill_1
XFILLER_10_1027 VPWR VGND sg13g2_fill_2
X_5445__110 VPWR VGND net110 sg13g2_tiehi
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_17_925 VPWR VGND sg13g2_decap_8
XFILLER_28_251 VPWR VGND sg13g2_fill_2
XFILLER_29_796 VPWR VGND sg13g2_fill_1
XFILLER_44_755 VPWR VGND sg13g2_fill_1
XFILLER_43_232 VPWR VGND sg13g2_decap_4
XFILLER_16_446 VPWR VGND sg13g2_decap_8
XFILLER_32_906 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_23_clk clknet_3_4__leaf_clk clknet_leaf_23_clk VPWR VGND sg13g2_buf_8
XFILLER_31_449 VPWR VGND sg13g2_fill_1
XFILLER_8_634 VPWR VGND sg13g2_fill_1
XFILLER_4_873 VPWR VGND sg13g2_decap_8
X_3180_ VGND VPWR _2280_ net682 _0032_ _0395_ sg13g2_a21oi_1
XFILLER_39_516 VPWR VGND sg13g2_decap_8
XFILLER_39_549 VPWR VGND sg13g2_fill_2
XFILLER_14_4 VPWR VGND sg13g2_fill_2
XFILLER_19_284 VPWR VGND sg13g2_fill_1
XFILLER_34_221 VPWR VGND sg13g2_decap_8
XFILLER_34_276 VPWR VGND sg13g2_fill_1
X_2964_ VGND VPWR _2190_ net691 _2318_ net789 sg13g2_a21oi_1
Xclkbuf_leaf_14_clk clknet_3_2__leaf_clk clknet_leaf_14_clk VPWR VGND sg13g2_buf_8
X_4703_ net819 VPWR _1650_ VGND net1088 net628 sg13g2_o21ai_1
XFILLER_31_961 VPWR VGND sg13g2_decap_8
XFILLER_33_1016 VPWR VGND sg13g2_decap_8
XFILLER_33_1027 VPWR VGND sg13g2_fill_2
X_2895_ net1166 _2249_ VPWR VGND sg13g2_inv_4
X_4634_ VPWR VGND net616 _1582_ _1547_ _1309_ _1583_ _1546_ sg13g2_a221oi_1
X_4565_ _1224_ _1304_ _1321_ _1515_ VPWR VGND sg13g2_nor3_1
X_3516_ _2249_ net586 _0689_ VPWR VGND sg13g2_nor2_1
X_4496_ _1074_ VPWR _1447_ VGND _1226_ _1314_ sg13g2_o21ai_1
X_3447_ _0623_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] net594 VPWR VGND sg13g2_nand2_1
X_3378_ _0556_ _0554_ _0555_ _2271_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] VPWR VGND
+ sg13g2_a22oi_1
XFILLER_40_1009 VPWR VGND sg13g2_decap_8
X_5117_ VGND VPWR net714 net747 _2056_ _1275_ sg13g2_a21oi_1
X_5048_ _1944_ _1954_ _1989_ VPWR VGND sg13g2_nor2_1
Xheichips25_tiny_wrapper_20 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_26_722 VPWR VGND sg13g2_fill_2
XFILLER_25_298 VPWR VGND sg13g2_fill_1
XFILLER_22_950 VPWR VGND sg13g2_decap_8
XFILLER_4_114 VPWR VGND sg13g2_fill_2
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_44_530 VPWR VGND sg13g2_fill_1
XFILLER_17_788 VPWR VGND sg13g2_fill_2
XFILLER_17_799 VPWR VGND sg13g2_fill_1
XFILLER_13_950 VPWR VGND sg13g2_decap_8
XFILLER_20_909 VPWR VGND sg13g2_decap_8
XFILLER_9_965 VPWR VGND sg13g2_decap_8
X_4350_ falu_i.falutop.alu_inst.op\[1\] falu_i.falutop.alu_inst.op\[0\] net771 _1303_
+ VPWR VGND sg13g2_nor3_2
X_3301_ VPWR VGND _0477_ _2255_ _0482_ _2257_ _0483_ _0478_ sg13g2_a221oi_1
X_4281_ _1231_ _1232_ _1234_ VPWR VGND sg13g2_nor2_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk clknet_leaf_3_clk VPWR VGND sg13g2_buf_8
X_3232_ _2270_ _2271_ _0427_ _0431_ VPWR VGND sg13g2_nor3_2
X_3163_ net811 VPWR _0387_ VGND ppwm_i.u_ppwm.pwm_value\[0\] net681 sg13g2_o21ai_1
X_3094_ net816 VPWR _2444_ VGND net848 _2443_ sg13g2_o21ai_1
XFILLER_22_213 VPWR VGND sg13g2_fill_1
XFILLER_23_758 VPWR VGND sg13g2_decap_8
XFILLER_10_408 VPWR VGND sg13g2_fill_1
XFILLER_11_909 VPWR VGND sg13g2_decap_8
X_3996_ net652 _1029_ _1030_ VPWR VGND sg13g2_nor2_2
X_2947_ net769 _2301_ VPWR VGND sg13g2_inv_4
X_4617_ _1566_ _1494_ _1565_ VPWR VGND sg13g2_xnor2_1
X_2878_ VPWR _2232_ net560 VGND sg13g2_inv_1
Xhold420 _0309_ VPWR VGND net1072 sg13g2_dlygate4sd3_1
Xhold442 ppwm_i.u_ppwm.u_pwm.counter\[8\] VPWR VGND net1094 sg13g2_dlygate4sd3_1
Xhold431 falu_i.falutop.i2c_inst.result\[4\] VPWR VGND net1083 sg13g2_dlygate4sd3_1
Xhold453 falu_i.falutop.data_in\[14\] VPWR VGND net1105 sg13g2_dlygate4sd3_1
X_4548_ _1497_ VPWR _1498_ VGND _1434_ _1495_ sg13g2_o21ai_1
Xhold486 _0320_ VPWR VGND net1138 sg13g2_dlygate4sd3_1
Xhold464 falu_i.falutop.div_inst.rem\[0\] VPWR VGND net1116 sg13g2_dlygate4sd3_1
X_4479_ _1428_ _1233_ _1430_ VPWR VGND sg13g2_xor2_1
Xhold475 falu_i.falutop.data_in\[2\] VPWR VGND net1127 sg13g2_dlygate4sd3_1
Xhold497 _0313_ VPWR VGND net1149 sg13g2_dlygate4sd3_1
XFILLER_38_24 VPWR VGND sg13g2_decap_4
XFILLER_18_508 VPWR VGND sg13g2_fill_1
XFILLER_46_839 VPWR VGND sg13g2_fill_2
XFILLER_45_327 VPWR VGND sg13g2_fill_1
XFILLER_14_703 VPWR VGND sg13g2_fill_1
XFILLER_14_747 VPWR VGND sg13g2_decap_4
XFILLER_16_1000 VPWR VGND sg13g2_decap_8
X_5488__305 VPWR VGND net305 sg13g2_tiehi
XFILLER_10_964 VPWR VGND sg13g2_decap_8
XFILLER_6_913 VPWR VGND sg13g2_decap_8
XFILLER_5_423 VPWR VGND sg13g2_fill_1
X_5306__88 VPWR VGND net88 sg13g2_tiehi
X_5421__208 VPWR VGND net208 sg13g2_tiehi
XFILLER_36_305 VPWR VGND sg13g2_fill_1
XFILLER_45_894 VPWR VGND sg13g2_decap_8
X_3850_ VGND VPWR _2204_ net664 _0144_ _0953_ sg13g2_a21oi_1
XFILLER_32_544 VPWR VGND sg13g2_fill_2
X_2801_ VPWR _2155_ net1051 VGND sg13g2_inv_1
X_3781_ net827 VPWR _0919_ VGND net504 net660 sg13g2_o21ai_1
X_5520_ net198 VGND VPWR _0279_ falu_i.falutop.div_inst.rem\[7\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_5451_ net82 VGND VPWR _0210_ ppwm_i.u_ppwm.u_mem.memory\[110\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_5382_ net288 VGND VPWR net970 ppwm_i.u_ppwm.u_mem.memory\[41\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_4402_ _1354_ _1350_ _1351_ VPWR VGND sg13g2_xnor2_1
X_4333_ VGND VPWR _1286_ net725 net721 sg13g2_or2_1
XFILLER_5_83 VPWR VGND sg13g2_fill_2
X_4264_ _1214_ _1216_ _1217_ VPWR VGND sg13g2_nor2_1
X_3215_ net809 VPWR _0420_ VGND _2273_ _0418_ sg13g2_o21ai_1
X_4195_ net803 VPWR _1168_ VGND net1119 net635 sg13g2_o21ai_1
X_3146_ VGND VPWR net802 _0374_ _0018_ _0375_ sg13g2_a21oi_1
XFILLER_39_198 VPWR VGND sg13g2_fill_2
X_3077_ _2429_ net1039 net821 VPWR VGND sg13g2_nand2_1
XFILLER_42_319 VPWR VGND sg13g2_decap_4
XFILLER_36_850 VPWR VGND sg13g2_decap_8
XFILLER_36_861 VPWR VGND sg13g2_fill_2
XFILLER_39_1022 VPWR VGND sg13g2_decap_8
XFILLER_35_360 VPWR VGND sg13g2_fill_1
XFILLER_35_371 VPWR VGND sg13g2_fill_1
XFILLER_11_717 VPWR VGND sg13g2_decap_4
X_3979_ net836 VPWR _1018_ VGND net461 net667 sg13g2_o21ai_1
XFILLER_3_938 VPWR VGND sg13g2_decap_8
XFILLER_2_437 VPWR VGND sg13g2_fill_1
Xhold261 _0093_ VPWR VGND net913 sg13g2_dlygate4sd3_1
Xhold250 _0229_ VPWR VGND net902 sg13g2_dlygate4sd3_1
Xhold272 ppwm_i.u_ppwm.u_pwm.cmp_value\[8\] VPWR VGND net924 sg13g2_dlygate4sd3_1
Xhold294 _0238_ VPWR VGND net946 sg13g2_dlygate4sd3_1
Xhold283 _1045_ VPWR VGND net935 sg13g2_dlygate4sd3_1
Xfanout730 falu_i.falutop.alu_data_in\[11\] net730 VPWR VGND sg13g2_buf_8
Xfanout741 net742 net741 VPWR VGND sg13g2_buf_8
X_5344__364 VPWR VGND net364 sg13g2_tiehi
Xfanout774 net775 net774 VPWR VGND sg13g2_buf_1
Xfanout752 net754 net752 VPWR VGND sg13g2_buf_8
Xfanout763 net764 net763 VPWR VGND sg13g2_buf_1
Xfanout785 net1196 net785 VPWR VGND sg13g2_buf_8
XFILLER_19_828 VPWR VGND sg13g2_decap_8
Xfanout796 net797 net796 VPWR VGND sg13g2_buf_8
XFILLER_42_820 VPWR VGND sg13g2_fill_1
XFILLER_14_500 VPWR VGND sg13g2_decap_4
XFILLER_42_853 VPWR VGND sg13g2_fill_2
XFILLER_26_393 VPWR VGND sg13g2_decap_4
XFILLER_10_761 VPWR VGND sg13g2_fill_2
XFILLER_6_732 VPWR VGND sg13g2_fill_1
XFILLER_5_297 VPWR VGND sg13g2_fill_1
XFILLER_2_960 VPWR VGND sg13g2_decap_8
XFILLER_49_441 VPWR VGND sg13g2_decap_8
X_3000_ ppwm_i.u_ppwm.u_mem.memory\[16\] net693 _2354_ VPWR VGND sg13g2_and2_1
XFILLER_49_496 VPWR VGND sg13g2_fill_2
XFILLER_36_124 VPWR VGND sg13g2_fill_2
X_5395__262 VPWR VGND net262 sg13g2_tiehi
XFILLER_18_872 VPWR VGND sg13g2_decap_8
X_4951_ _1854_ VPWR _1894_ VGND _1853_ _1855_ sg13g2_o21ai_1
XFILLER_17_360 VPWR VGND sg13g2_fill_2
X_3902_ VGND VPWR _2185_ net671 _0170_ _0979_ sg13g2_a21oi_1
X_4882_ _1827_ _1789_ _1826_ VPWR VGND sg13g2_nand2_1
XFILLER_32_330 VPWR VGND sg13g2_fill_2
X_3833_ net830 VPWR _0945_ VGND net481 net664 sg13g2_o21ai_1
X_3764_ VGND VPWR _2234_ net644 _0101_ _0910_ sg13g2_a21oi_1
X_3695_ _0856_ _2238_ net600 VPWR VGND sg13g2_xnor2_1
XFILLER_9_581 VPWR VGND sg13g2_decap_8
X_5503_ net269 VGND VPWR net1055 falu_i.falutop.div_inst.b1\[7\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
X_5434_ net155 VGND VPWR _0193_ ppwm_i.u_ppwm.u_mem.memory\[93\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_5365_ net322 VGND VPWR _0124_ ppwm_i.u_ppwm.u_mem.memory\[24\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_4316_ _1268_ _1264_ _1225_ _1269_ VPWR VGND sg13g2_a21o_1
X_5296_ net105 VGND VPWR _0058_ ppwm_i.u_ppwm.global_counter\[13\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_4247_ _1207_ net489 _1105_ VPWR VGND sg13g2_nand2_1
X_4178_ _1154_ net479 net568 VPWR VGND sg13g2_nand2_1
X_3129_ net820 VPWR _0364_ VGND net899 _0363_ sg13g2_o21ai_1
XFILLER_27_146 VPWR VGND sg13g2_fill_2
XFILLER_27_157 VPWR VGND sg13g2_fill_1
XFILLER_36_680 VPWR VGND sg13g2_fill_2
XFILLER_35_69 VPWR VGND sg13g2_fill_2
XFILLER_24_886 VPWR VGND sg13g2_decap_8
XFILLER_11_536 VPWR VGND sg13g2_decap_4
XFILLER_23_396 VPWR VGND sg13g2_decap_4
XFILLER_46_400 VPWR VGND sg13g2_decap_8
Xfanout582 net583 net582 VPWR VGND sg13g2_buf_8
Xfanout571 _0628_ net571 VPWR VGND sg13g2_buf_8
Xfanout593 net597 net593 VPWR VGND sg13g2_buf_8
XFILLER_47_967 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_fill_1
XFILLER_20_1007 VPWR VGND sg13g2_decap_8
X_5460__46 VPWR VGND net46 sg13g2_tiehi
XFILLER_14_374 VPWR VGND sg13g2_fill_2
XFILLER_15_875 VPWR VGND sg13g2_decap_8
XFILLER_6_562 VPWR VGND sg13g2_decap_8
X_3480_ VPWR _0655_ _0654_ VGND sg13g2_inv_1
XFILLER_6_584 VPWR VGND sg13g2_decap_4
X_5150_ VGND VPWR net638 _2087_ _2088_ net630 sg13g2_a21oi_1
X_5081_ _2021_ _1944_ _1987_ VPWR VGND sg13g2_nand2_2
X_4101_ _1104_ net778 _1101_ VPWR VGND sg13g2_nand2_2
X_4032_ _1058_ _2442_ _0901_ VPWR VGND sg13g2_nand2_1
XFILLER_38_967 VPWR VGND sg13g2_decap_8
XFILLER_37_444 VPWR VGND sg13g2_fill_1
X_4934_ _1878_ _1841_ _1876_ VPWR VGND sg13g2_nand2b_1
XFILLER_21_812 VPWR VGND sg13g2_decap_8
XFILLER_36_1025 VPWR VGND sg13g2_decap_4
X_4865_ net718 net761 net723 _1810_ VPWR VGND net755 sg13g2_nand4_1
X_4796_ net746 net706 _1742_ VPWR VGND sg13g2_nor2_1
XFILLER_21_889 VPWR VGND sg13g2_decap_8
X_3816_ VGND VPWR _2215_ net654 _0127_ _0936_ sg13g2_a21oi_1
X_3747_ falu_i.falutop.i2c_inst.data_in\[16\] net686 _0903_ VPWR VGND sg13g2_nor2_1
X_3678_ _0841_ _0840_ _0839_ VPWR VGND sg13g2_nand2b_1
X_5417_ net218 VGND VPWR _0176_ ppwm_i.u_ppwm.u_mem.memory\[76\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_5348_ net356 VGND VPWR _0107_ ppwm_i.u_ppwm.u_mem.memory\[7\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_5279_ net138 VGND VPWR _0041_ ppwm_i.u_ppwm.u_pwm.counter\[7\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_2
X_5263__170 VPWR VGND net170 sg13g2_tiehi
XFILLER_29_956 VPWR VGND sg13g2_decap_8
XFILLER_44_937 VPWR VGND sg13g2_decap_8
XFILLER_12_801 VPWR VGND sg13g2_fill_1
XFILLER_24_650 VPWR VGND sg13g2_decap_8
XFILLER_11_322 VPWR VGND sg13g2_fill_2
XFILLER_24_683 VPWR VGND sg13g2_decap_8
XFILLER_12_867 VPWR VGND sg13g2_decap_8
XFILLER_7_29 VPWR VGND sg13g2_fill_2
XFILLER_3_521 VPWR VGND sg13g2_fill_2
XFILLER_3_543 VPWR VGND sg13g2_fill_1
XFILLER_19_400 VPWR VGND sg13g2_fill_1
X_2980_ _2332_ _2333_ _2331_ _2334_ VPWR VGND sg13g2_nand3_1
XFILLER_14_160 VPWR VGND sg13g2_decap_8
XFILLER_15_694 VPWR VGND sg13g2_decap_4
X_4650_ _1536_ _1597_ _1598_ VPWR VGND sg13g2_nor2_1
X_3601_ net584 _0677_ _0770_ VPWR VGND sg13g2_nor2_1
XFILLER_7_860 VPWR VGND sg13g2_decap_8
X_4581_ net717 net754 net736 _1530_ VPWR VGND sg13g2_nand3_1
X_3532_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] _0704_ net588 _0705_ VPWR VGND sg13g2_mux2_1
XFILLER_6_392 VPWR VGND sg13g2_decap_8
XFILLER_6_381 VPWR VGND sg13g2_fill_1
X_3463_ net594 ppwm_i.u_ppwm.global_counter\[0\] _0639_ VPWR VGND sg13g2_nor2b_1
X_5202_ _2118_ falu_i.falutop.data_in\[3\] _2117_ VPWR VGND sg13g2_xnor2_1
X_5133_ _2072_ net773 _2047_ VPWR VGND sg13g2_nand2_1
X_3394_ _0571_ VPWR _0572_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] _2266_ sg13g2_o21ai_1
XFILLER_35_0 VPWR VGND sg13g2_decap_4
X_5064_ _2004_ _1984_ _2005_ VPWR VGND sg13g2_nor2b_1
X_4015_ ppwm_i.u_ppwm.u_mem.bit_count\[4\] _0397_ _1034_ _1044_ VPWR VGND sg13g2_nor3_1
XFILLER_26_937 VPWR VGND sg13g2_decap_8
XFILLER_25_447 VPWR VGND sg13g2_fill_1
X_4917_ _1752_ _1858_ _1859_ _1861_ VPWR VGND sg13g2_or3_1
X_4848_ net742 net706 _1793_ VPWR VGND sg13g2_nor2_1
X_4779_ _1310_ _1724_ _1725_ VPWR VGND sg13g2_nor2_1
XFILLER_10_1006 VPWR VGND sg13g2_decap_8
XFILLER_0_546 VPWR VGND sg13g2_fill_2
XFILLER_17_904 VPWR VGND sg13g2_decap_8
XFILLER_25_981 VPWR VGND sg13g2_decap_8
X_5569__72 VPWR VGND net72 sg13g2_tiehi
XFILLER_40_995 VPWR VGND sg13g2_decap_8
XFILLER_8_646 VPWR VGND sg13g2_decap_4
XFILLER_12_697 VPWR VGND sg13g2_fill_1
XFILLER_11_196 VPWR VGND sg13g2_decap_8
XFILLER_4_852 VPWR VGND sg13g2_decap_8
XFILLER_35_745 VPWR VGND sg13g2_fill_1
XFILLER_34_255 VPWR VGND sg13g2_fill_2
X_2963_ ppwm_i.u_ppwm.u_mem.memory\[57\] _2310_ _2317_ VPWR VGND sg13g2_nor2_1
X_4702_ _1648_ _1649_ _0300_ VPWR VGND sg13g2_nor2_1
XFILLER_31_940 VPWR VGND sg13g2_decap_8
X_2894_ ppwm_i.u_ppwm.pwm_value\[4\] _2248_ VPWR VGND sg13g2_inv_4
X_4633_ _1579_ _1581_ _1569_ _1582_ VPWR VGND sg13g2_nand3_1
XFILLER_30_494 VPWR VGND sg13g2_fill_2
X_4564_ _1514_ _1224_ _1319_ VPWR VGND sg13g2_nand2_1
X_3515_ _0670_ VPWR _0688_ VGND _2250_ net586 sg13g2_o21ai_1
X_4495_ _1441_ VPWR _1446_ VGND _1374_ _1444_ sg13g2_o21ai_1
X_5284__129 VPWR VGND net129 sg13g2_tiehi
X_3446_ _2375_ _0621_ _0622_ VPWR VGND sg13g2_nor2_2
X_3377_ _0555_ ppwm_i.u_ppwm.global_counter\[1\] _2242_ ppwm_i.u_ppwm.global_counter\[2\]
+ _2241_ VPWR VGND sg13g2_a22oi_1
X_5116_ _2021_ VPWR _2055_ VGND _2023_ _2032_ sg13g2_o21ai_1
X_5047_ _1988_ _1947_ _1987_ VPWR VGND sg13g2_xnor2_1
Xheichips25_tiny_wrapper_21 VPWR VGND uio_out[5] sg13g2_tielo
Xheichips25_tiny_wrapper_10 VPWR VGND uio_oe[2] sg13g2_tielo
XFILLER_14_929 VPWR VGND sg13g2_decap_8
X_5949_ falu_i.falutop.i2c_inst.sda_o net6 VPWR VGND sg13g2_buf_2
XFILLER_40_269 VPWR VGND sg13g2_fill_1
XFILLER_5_638 VPWR VGND sg13g2_decap_8
XFILLER_49_1013 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_fill_2
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_49_815 VPWR VGND sg13g2_decap_4
XFILLER_49_859 VPWR VGND sg13g2_decap_8
XFILLER_48_369 VPWR VGND sg13g2_fill_1
XFILLER_1_1015 VPWR VGND sg13g2_decap_8
XFILLER_17_745 VPWR VGND sg13g2_fill_2
X_5354__344 VPWR VGND net344 sg13g2_tiehi
XFILLER_31_214 VPWR VGND sg13g2_fill_1
XFILLER_9_944 VPWR VGND sg13g2_decap_8
XFILLER_12_461 VPWR VGND sg13g2_fill_2
XFILLER_8_487 VPWR VGND sg13g2_fill_1
X_3300_ _2330_ _0478_ _0482_ VPWR VGND sg13g2_nor2_2
XFILLER_4_682 VPWR VGND sg13g2_decap_8
X_4280_ _1233_ net741 net766 VPWR VGND sg13g2_nand2_2
XFILLER_3_192 VPWR VGND sg13g2_fill_2
X_3231_ net795 _0429_ _0430_ _0048_ VPWR VGND sg13g2_nor3_1
X_3162_ _2274_ _0384_ _2273_ _0386_ VPWR VGND _0385_ sg13g2_nand4_1
X_3093_ net1014 _2439_ _2443_ VPWR VGND sg13g2_nor2_1
XFILLER_23_737 VPWR VGND sg13g2_decap_8
X_3995_ _1029_ net1051 _1025_ VPWR VGND sg13g2_nand2_1
X_2946_ _2300_ net771 VPWR VGND sg13g2_inv_2
X_2877_ VPWR _2231_ net483 VGND sg13g2_inv_1
X_4616_ _1565_ _1548_ _1562_ VPWR VGND sg13g2_xnor2_1
Xhold410 falu_i.falutop.i2c_inst.result\[10\] VPWR VGND net1062 sg13g2_dlygate4sd3_1
Xhold443 _0042_ VPWR VGND net1095 sg13g2_dlygate4sd3_1
Xhold454 falu_i.falutop.div_inst.rem\[5\] VPWR VGND net1106 sg13g2_dlygate4sd3_1
Xhold432 falu_i.falutop.i2c_inst.result\[5\] VPWR VGND net1084 sg13g2_dlygate4sd3_1
XFILLER_2_608 VPWR VGND sg13g2_fill_2
Xhold421 falu_i.falutop.data_in\[6\] VPWR VGND net1073 sg13g2_dlygate4sd3_1
X_4547_ _1318_ _1496_ _1497_ VPWR VGND sg13g2_nor2_1
Xhold487 ppwm_i.u_ppwm.global_counter\[9\] VPWR VGND net1139 sg13g2_dlygate4sd3_1
X_4478_ _1233_ _1428_ _1429_ VPWR VGND sg13g2_nor2_1
Xhold476 _0315_ VPWR VGND net1128 sg13g2_dlygate4sd3_1
Xhold465 ppwm_i.u_ppwm.u_pwm.counter\[1\] VPWR VGND net1117 sg13g2_dlygate4sd3_1
X_3429_ _2361_ _2375_ net419 _0606_ VPWR VGND net582 sg13g2_nand4_1
Xhold498 falu_i.falutop.i2c_inst.counter\[4\] VPWR VGND net1150 sg13g2_dlygate4sd3_1
XFILLER_38_47 VPWR VGND sg13g2_fill_2
XFILLER_38_380 VPWR VGND sg13g2_fill_1
XFILLER_13_214 VPWR VGND sg13g2_decap_4
XFILLER_10_943 VPWR VGND sg13g2_decap_8
XFILLER_6_969 VPWR VGND sg13g2_decap_8
X_5321__59 VPWR VGND net59 sg13g2_tiehi
XFILLER_0_195 VPWR VGND sg13g2_decap_8
XFILLER_0_184 VPWR VGND sg13g2_fill_2
XFILLER_0_173 VPWR VGND sg13g2_fill_2
XFILLER_48_155 VPWR VGND sg13g2_fill_1
XFILLER_17_553 VPWR VGND sg13g2_fill_1
X_5471__343 VPWR VGND net343 sg13g2_tiehi
X_2800_ _2154_ net1006 VPWR VGND sg13g2_inv_2
X_3780_ VGND VPWR _2228_ net662 _0109_ _0918_ sg13g2_a21oi_1
XFILLER_9_741 VPWR VGND sg13g2_decap_8
XFILLER_12_280 VPWR VGND sg13g2_fill_1
XFILLER_8_251 VPWR VGND sg13g2_fill_1
XFILLER_8_240 VPWR VGND sg13g2_decap_8
X_5450_ net86 VGND VPWR _0209_ ppwm_i.u_ppwm.u_mem.memory\[109\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_4401_ _1353_ _1350_ _1352_ VPWR VGND sg13g2_nand2_1
X_5381_ net290 VGND VPWR net456 ppwm_i.u_ppwm.u_mem.memory\[40\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_4332_ net730 net736 _1285_ VPWR VGND sg13g2_nor2_1
XFILLER_4_490 VPWR VGND sg13g2_fill_1
X_4263_ net722 net750 _1216_ VPWR VGND sg13g2_nor2_2
X_3214_ VGND VPWR _2274_ _0417_ _0042_ _0419_ sg13g2_a21oi_1
X_4194_ _1166_ VPWR _1167_ VGND net494 net568 sg13g2_o21ai_1
X_3145_ net804 VPWR _0375_ VGND net861 _0374_ sg13g2_o21ai_1
X_3076_ net980 net385 _2428_ VPWR VGND sg13g2_nor2_1
XFILLER_39_1001 VPWR VGND sg13g2_decap_8
X_3978_ VGND VPWR _2158_ net667 _0208_ _1017_ sg13g2_a21oi_1
X_2929_ VPWR _2283_ net426 VGND sg13g2_inv_1
XFILLER_40_37 VPWR VGND sg13g2_fill_2
X_5579_ net263 VGND VPWR net476 falu_i.falutop.div_inst.a\[2\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
XFILLER_3_917 VPWR VGND sg13g2_decap_8
Xhold251 ppwm_i.u_ppwm.u_mem.memory\[66\] VPWR VGND net903 sg13g2_dlygate4sd3_1
Xhold240 _0331_ VPWR VGND net892 sg13g2_dlygate4sd3_1
Xhold262 ppwm_i.u_ppwm.u_mem.memory\[105\] VPWR VGND net914 sg13g2_dlygate4sd3_1
Xhold273 _0032_ VPWR VGND net925 sg13g2_dlygate4sd3_1
Xhold295 falu_i.falutop.div_inst.val\[3\] VPWR VGND net947 sg13g2_dlygate4sd3_1
Xhold284 _0219_ VPWR VGND net936 sg13g2_dlygate4sd3_1
XFILLER_49_79 VPWR VGND sg13g2_fill_2
Xfanout720 falu_i.falutop.alu_data_in\[14\] net720 VPWR VGND sg13g2_buf_8
Xfanout731 falu_i.falutop.alu_data_in\[11\] net731 VPWR VGND sg13g2_buf_8
Xfanout742 falu_i.falutop.alu_data_in\[9\] net742 VPWR VGND sg13g2_buf_8
Xfanout753 net754 net753 VPWR VGND sg13g2_buf_1
Xfanout775 net776 net775 VPWR VGND sg13g2_buf_1
Xfanout764 net765 net764 VPWR VGND sg13g2_buf_2
Xfanout786 net1192 net786 VPWR VGND sg13g2_buf_8
Xfanout797 _2294_ net797 VPWR VGND sg13g2_buf_8
XFILLER_45_125 VPWR VGND sg13g2_decap_8
XFILLER_42_810 VPWR VGND sg13g2_fill_1
XFILLER_14_545 VPWR VGND sg13g2_decap_8
XFILLER_41_353 VPWR VGND sg13g2_fill_1
X_5273__150 VPWR VGND net150 sg13g2_tiehi
XFILLER_14_71 VPWR VGND sg13g2_decap_8
XFILLER_6_711 VPWR VGND sg13g2_decap_8
XFILLER_49_420 VPWR VGND sg13g2_decap_8
XFILLER_7_1021 VPWR VGND sg13g2_decap_8
XFILLER_1_493 VPWR VGND sg13g2_fill_2
XFILLER_49_475 VPWR VGND sg13g2_decap_8
XFILLER_18_851 VPWR VGND sg13g2_decap_8
X_4950_ _1868_ VPWR _1893_ VGND _1851_ _1869_ sg13g2_o21ai_1
X_3901_ net834 VPWR _0979_ VGND ppwm_i.u_ppwm.u_mem.memory\[70\] net669 sg13g2_o21ai_1
X_4881_ _1825_ _1747_ _1826_ VPWR VGND sg13g2_xor2_1
XFILLER_33_843 VPWR VGND sg13g2_decap_4
X_3832_ VGND VPWR _2210_ net642 _0135_ _0944_ sg13g2_a21oi_1
XFILLER_33_898 VPWR VGND sg13g2_fill_1
X_5502_ net271 VGND VPWR _0261_ falu_i.falutop.div_inst.b1\[6\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_2
X_3763_ net827 VPWR _0910_ VGND ppwm_i.u_ppwm.u_mem.memory\[2\] net644 sg13g2_o21ai_1
X_3694_ VPWR VGND _0855_ net795 _0852_ _2239_ _0086_ net569 sg13g2_a221oi_1
X_5433_ net159 VGND VPWR _0192_ ppwm_i.u_ppwm.u_mem.memory\[92\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_5364_ net324 VGND VPWR net403 ppwm_i.u_ppwm.u_mem.memory\[23\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_4315_ VGND VPWR _1268_ _1267_ _1229_ sg13g2_or2_1
X_5295_ net107 VGND VPWR _0057_ ppwm_i.u_ppwm.global_counter\[12\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_4246_ _1206_ VPWR _0287_ VGND _1098_ _1155_ sg13g2_o21ai_1
X_4177_ VGND VPWR _2146_ net636 _0271_ _1153_ sg13g2_a21oi_1
X_3128_ _2446_ _0360_ _0363_ VPWR VGND sg13g2_nor2_1
XFILLER_28_648 VPWR VGND sg13g2_fill_2
X_3059_ _2413_ net696 _2212_ net700 _2198_ VPWR VGND sg13g2_a22oi_1
XFILLER_43_618 VPWR VGND sg13g2_fill_2
XFILLER_24_865 VPWR VGND sg13g2_decap_8
XFILLER_35_191 VPWR VGND sg13g2_decap_8
Xfanout583 _0530_ net583 VPWR VGND sg13g2_buf_8
XFILLER_19_604 VPWR VGND sg13g2_decap_4
Xfanout572 net573 net572 VPWR VGND sg13g2_buf_8
XFILLER_47_946 VPWR VGND sg13g2_decap_8
Xfanout594 net596 net594 VPWR VGND sg13g2_buf_8
XFILLER_14_331 VPWR VGND sg13g2_decap_8
XFILLER_15_854 VPWR VGND sg13g2_decap_8
XFILLER_41_161 VPWR VGND sg13g2_decap_4
XFILLER_2_780 VPWR VGND sg13g2_decap_8
X_5080_ _1990_ _1999_ _2020_ VPWR VGND sg13g2_nor2_1
X_4100_ net778 _1101_ _1103_ VPWR VGND sg13g2_and2_1
X_4031_ net459 net1015 _1057_ VPWR VGND sg13g2_nor2_1
XFILLER_49_283 VPWR VGND sg13g2_decap_8
XFILLER_38_946 VPWR VGND sg13g2_decap_8
XFILLER_37_401 VPWR VGND sg13g2_decap_8
XFILLER_25_629 VPWR VGND sg13g2_decap_8
X_4933_ _1841_ _1876_ _1877_ VPWR VGND sg13g2_nor2b_1
XFILLER_36_1004 VPWR VGND sg13g2_decap_8
X_4864_ net723 net718 net761 net755 _1809_ VPWR VGND sg13g2_and4_1
X_4795_ _1689_ VPWR _1741_ VGND _1687_ _1690_ sg13g2_o21ai_1
XFILLER_21_868 VPWR VGND sg13g2_decap_8
X_3815_ net824 VPWR _0936_ VGND ppwm_i.u_ppwm.u_mem.memory\[27\] net654 sg13g2_o21ai_1
X_3746_ falu_i.falutop.i2c_inst.state\[0\] net804 net459 _0902_ VPWR VGND sg13g2_nand3_1
X_5416_ net220 VGND VPWR _0175_ ppwm_i.u_ppwm.u_mem.memory\[75\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_3677_ _0840_ _2240_ net586 VPWR VGND sg13g2_nand2_1
XFILLER_0_706 VPWR VGND sg13g2_decap_4
X_5347_ net358 VGND VPWR _0106_ ppwm_i.u_ppwm.u_mem.memory\[6\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_5278_ net140 VGND VPWR net1068 ppwm_i.u_ppwm.u_pwm.counter\[6\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_1
XFILLER_47_209 VPWR VGND sg13g2_fill_2
X_4229_ net781 _2149_ _1194_ VPWR VGND sg13g2_nor2_1
XFILLER_29_935 VPWR VGND sg13g2_decap_8
XFILLER_44_916 VPWR VGND sg13g2_decap_8
X_5294__109 VPWR VGND net109 sg13g2_tiehi
XFILLER_11_312 VPWR VGND sg13g2_fill_1
XFILLER_12_846 VPWR VGND sg13g2_decap_8
XFILLER_8_817 VPWR VGND sg13g2_decap_4
XFILLER_23_194 VPWR VGND sg13g2_decap_8
XFILLER_8_839 VPWR VGND sg13g2_decap_8
X_5526__169 VPWR VGND net169 sg13g2_tiehi
X_5242__211 VPWR VGND net211 sg13g2_tiehi
XFILLER_4_1013 VPWR VGND sg13g2_decap_8
XFILLER_47_743 VPWR VGND sg13g2_fill_1
XFILLER_19_456 VPWR VGND sg13g2_decap_8
XFILLER_35_949 VPWR VGND sg13g2_decap_8
XFILLER_36_91 VPWR VGND sg13g2_fill_2
XFILLER_43_982 VPWR VGND sg13g2_decap_8
XFILLER_14_150 VPWR VGND sg13g2_decap_4
X_3600_ _0767_ _0768_ net575 _0769_ VPWR VGND sg13g2_nand3_1
X_4580_ _1529_ net737 net752 VPWR VGND sg13g2_nand2_1
X_3531_ _0703_ VPWR _0704_ VGND _2271_ net593 sg13g2_o21ai_1
X_5364__324 VPWR VGND net324 sg13g2_tiehi
X_3462_ _2419_ _0637_ _0638_ VPWR VGND sg13g2_nor2_1
X_5201_ _2096_ net777 _2117_ VPWR VGND sg13g2_nor2b_1
X_3393_ ppwm_i.u_ppwm.global_counter\[10\] ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] _0571_
+ VPWR VGND sg13g2_nor2b_1
X_5132_ _1590_ VPWR _2071_ VGND _2067_ _2070_ sg13g2_o21ai_1
X_5063_ _2003_ _1985_ _2004_ VPWR VGND sg13g2_xor2_1
XFILLER_37_231 VPWR VGND sg13g2_decap_8
X_4014_ net513 VPWR _0218_ VGND _1036_ _1043_ sg13g2_o21ai_1
XFILLER_38_787 VPWR VGND sg13g2_fill_2
XFILLER_26_916 VPWR VGND sg13g2_decap_8
Xheichips25_tiny_wrapper_8 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_40_429 VPWR VGND sg13g2_fill_2
X_4916_ _1752_ VPWR _1860_ VGND _1858_ _1859_ sg13g2_o21ai_1
XFILLER_33_470 VPWR VGND sg13g2_fill_2
X_4847_ _1754_ VPWR _1792_ VGND _1750_ _1755_ sg13g2_o21ai_1
XFILLER_21_654 VPWR VGND sg13g2_fill_2
X_4778_ _1660_ _1663_ _1722_ _1724_ VPWR VGND sg13g2_nor3_1
X_3729_ _0887_ _0884_ _0886_ VPWR VGND sg13g2_nand2_1
XFILLER_0_525 VPWR VGND sg13g2_fill_2
XFILLER_29_721 VPWR VGND sg13g2_fill_1
XFILLER_29_743 VPWR VGND sg13g2_decap_4
XFILLER_28_275 VPWR VGND sg13g2_decap_8
XFILLER_29_776 VPWR VGND sg13g2_fill_2
XFILLER_29_787 VPWR VGND sg13g2_decap_8
XFILLER_19_1010 VPWR VGND sg13g2_decap_8
XFILLER_25_960 VPWR VGND sg13g2_decap_8
XFILLER_43_289 VPWR VGND sg13g2_fill_1
XFILLER_31_418 VPWR VGND sg13g2_fill_1
XFILLER_40_974 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_decap_4
X_5336__32 VPWR VGND net32 sg13g2_tiehi
XFILLER_4_831 VPWR VGND sg13g2_decap_8
XFILLER_3_396 VPWR VGND sg13g2_fill_1
XFILLER_26_1014 VPWR VGND sg13g2_decap_8
XFILLER_19_231 VPWR VGND sg13g2_fill_1
XFILLER_47_90 VPWR VGND sg13g2_fill_2
XFILLER_19_242 VPWR VGND sg13g2_fill_2
XFILLER_23_919 VPWR VGND sg13g2_decap_8
XFILLER_16_993 VPWR VGND sg13g2_decap_8
X_2962_ _2314_ _2315_ _2316_ VPWR VGND sg13g2_and2_1
X_4701_ net819 VPWR _1649_ VGND net1084 net628 sg13g2_o21ai_1
X_5550__251 VPWR VGND net251 sg13g2_tiehi
X_2893_ net1188 _2247_ VPWR VGND sg13g2_inv_4
XFILLER_8_51 VPWR VGND sg13g2_fill_2
X_4632_ _1306_ _1580_ _1270_ _1581_ VPWR VGND sg13g2_nand3_1
XFILLER_30_451 VPWR VGND sg13g2_fill_1
XFILLER_31_996 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_4
X_4563_ _1289_ _1302_ net771 _1513_ VPWR VGND _1333_ sg13g2_nand4_1
XFILLER_7_680 VPWR VGND sg13g2_fill_2
X_4494_ _1445_ _1229_ _1383_ VPWR VGND sg13g2_nand2_1
X_3514_ net798 _0687_ _0074_ VPWR VGND sg13g2_nor2_1
X_3445_ _0621_ _2419_ _0620_ VPWR VGND sg13g2_nand2b_1
X_5481__323 VPWR VGND net323 sg13g2_tiehi
X_3376_ _0553_ VPWR _0554_ VGND _2242_ ppwm_i.u_ppwm.global_counter\[1\] sg13g2_o21ai_1
X_5115_ VGND VPWR _1994_ _2031_ _2054_ _2030_ sg13g2_a21oi_1
X_5046_ _1987_ _1652_ _1950_ VPWR VGND sg13g2_xnor2_1
Xheichips25_tiny_wrapper_22 VPWR VGND uio_out[6] sg13g2_tielo
Xheichips25_tiny_wrapper_11 VPWR VGND uio_oe[3] sg13g2_tielo
XFILLER_38_595 VPWR VGND sg13g2_fill_2
XFILLER_14_908 VPWR VGND sg13g2_decap_8
XFILLER_22_985 VPWR VGND sg13g2_decap_8
X_5318__65 VPWR VGND net65 sg13g2_tiehi
X_5562__133 VPWR VGND net133 sg13g2_tiehi
X_5333__35 VPWR VGND net35 sg13g2_tiehi
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_0_355 VPWR VGND sg13g2_decap_4
XFILLER_0_377 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_44_510 VPWR VGND sg13g2_decap_8
XFILLER_17_735 VPWR VGND sg13g2_decap_4
XFILLER_29_595 VPWR VGND sg13g2_fill_2
XFILLER_17_757 VPWR VGND sg13g2_fill_2
XFILLER_17_779 VPWR VGND sg13g2_fill_1
XFILLER_44_576 VPWR VGND sg13g2_decap_4
XFILLER_31_248 VPWR VGND sg13g2_fill_1
XFILLER_9_923 VPWR VGND sg13g2_decap_8
XFILLER_12_440 VPWR VGND sg13g2_fill_2
XFILLER_13_985 VPWR VGND sg13g2_decap_8
XFILLER_40_793 VPWR VGND sg13g2_decap_8
XFILLER_12_495 VPWR VGND sg13g2_fill_1
X_5580__255 VPWR VGND net255 sg13g2_tiehi
X_3230_ _2271_ _0427_ _0430_ VPWR VGND sg13g2_nor2_1
X_3161_ ppwm_i.u_ppwm.u_pwm.counter\[7\] ppwm_i.u_ppwm.u_pwm.counter\[6\] ppwm_i.u_ppwm.u_pwm.counter\[5\]
+ ppwm_i.u_ppwm.u_pwm.counter\[4\] _0385_ VPWR VGND sg13g2_nor4_1
X_3092_ _2442_ _2438_ _2437_ VPWR VGND sg13g2_nand2b_1
XFILLER_48_893 VPWR VGND sg13g2_decap_8
XFILLER_47_381 VPWR VGND sg13g2_fill_2
XFILLER_35_543 VPWR VGND sg13g2_fill_1
XFILLER_35_598 VPWR VGND sg13g2_fill_1
X_3994_ VGND VPWR net1051 _1021_ _1028_ net680 sg13g2_a21oi_1
X_2945_ _2299_ net772 VPWR VGND sg13g2_inv_2
X_2876_ VPWR _2230_ net451 VGND sg13g2_inv_1
X_4615_ _1548_ _1562_ _1564_ VPWR VGND sg13g2_nor2b_1
Xhold411 _0305_ VPWR VGND net1063 sg13g2_dlygate4sd3_1
X_4546_ _1434_ _1495_ _1496_ VPWR VGND sg13g2_and2_1
Xhold400 _1028_ VPWR VGND net1052 sg13g2_dlygate4sd3_1
Xhold433 falu_i.falutop.div_inst.b1\[5\] VPWR VGND net1085 sg13g2_dlygate4sd3_1
Xhold422 _2100_ VPWR VGND net1074 sg13g2_dlygate4sd3_1
Xhold444 ppwm_i.u_ppwm.global_counter\[0\] VPWR VGND net1096 sg13g2_dlygate4sd3_1
Xhold455 ppwm_i.u_ppwm.global_counter\[4\] VPWR VGND net1107 sg13g2_dlygate4sd3_1
X_4477_ _1428_ net745 net763 VPWR VGND sg13g2_nand2_1
Xhold466 _0403_ VPWR VGND net1118 sg13g2_dlygate4sd3_1
Xhold477 ppwm_i.u_ppwm.global_counter\[13\] VPWR VGND net1129 sg13g2_dlygate4sd3_1
Xhold488 _0441_ VPWR VGND net1140 sg13g2_dlygate4sd3_1
X_3428_ net821 _0605_ _0070_ VPWR VGND sg13g2_and2_1
Xhold499 ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] VPWR VGND net1151 sg13g2_dlygate4sd3_1
X_3359_ _0537_ _0535_ _0536_ ppwm_i.u_ppwm.global_counter\[2\] _2250_ VPWR VGND sg13g2_a22oi_1
X_5557__202 VPWR VGND net202 sg13g2_tiehi
XFILLER_45_307 VPWR VGND sg13g2_fill_2
XFILLER_39_860 VPWR VGND sg13g2_decap_4
X_5029_ _1834_ VPWR _1971_ VGND _1282_ _1970_ sg13g2_o21ai_1
XFILLER_26_521 VPWR VGND sg13g2_decap_4
XFILLER_38_392 VPWR VGND sg13g2_decap_8
XFILLER_14_738 VPWR VGND sg13g2_decap_4
XFILLER_10_922 VPWR VGND sg13g2_decap_8
XFILLER_22_782 VPWR VGND sg13g2_decap_8
XFILLER_6_948 VPWR VGND sg13g2_decap_8
XFILLER_10_999 VPWR VGND sg13g2_decap_8
XFILLER_49_602 VPWR VGND sg13g2_fill_2
XFILLER_0_152 VPWR VGND sg13g2_decap_8
XFILLER_23_1017 VPWR VGND sg13g2_decap_8
XFILLER_23_1028 VPWR VGND sg13g2_fill_1
XFILLER_49_668 VPWR VGND sg13g2_decap_8
XFILLER_44_373 VPWR VGND sg13g2_fill_2
XFILLER_17_576 VPWR VGND sg13g2_decap_4
XFILLER_32_502 VPWR VGND sg13g2_fill_1
XFILLER_9_764 VPWR VGND sg13g2_fill_2
X_4400_ VPWR _1352_ _1351_ VGND sg13g2_inv_1
X_5380_ net292 VGND VPWR _0139_ ppwm_i.u_ppwm.u_mem.memory\[39\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_5250__195 VPWR VGND net195 sg13g2_tiehi
X_4331_ net716 net710 _1284_ VPWR VGND sg13g2_nor2_2
X_4262_ _1215_ net724 net751 VPWR VGND sg13g2_nand2_2
X_3213_ _0419_ net809 _0418_ VPWR VGND sg13g2_nand2_1
X_4193_ _1166_ net568 _1165_ VPWR VGND sg13g2_nand2_1
XFILLER_39_156 VPWR VGND sg13g2_fill_1
X_3144_ _0344_ net1007 _0374_ VPWR VGND sg13g2_nor2_1
X_3075_ _2427_ _2308_ _2423_ VPWR VGND sg13g2_nand2_1
XFILLER_23_502 VPWR VGND sg13g2_fill_1
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_35_384 VPWR VGND sg13g2_fill_1
XFILLER_35_395 VPWR VGND sg13g2_decap_8
X_3977_ net838 VPWR _1017_ VGND ppwm_i.u_ppwm.u_mem.memory\[108\] net667 sg13g2_o21ai_1
X_2928_ VPWR _2282_ net492 VGND sg13g2_inv_1
X_2859_ VPWR _2213_ net516 VGND sg13g2_inv_1
X_5578_ net289 VGND VPWR net389 falu_i.falutop.div_inst.a\[1\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
Xhold241 ppwm_i.u_ppwm.u_mem.memory\[45\] VPWR VGND net893 sg13g2_dlygate4sd3_1
Xhold252 ppwm_i.u_ppwm.u_mem.memory\[68\] VPWR VGND net904 sg13g2_dlygate4sd3_1
XFILLER_2_428 VPWR VGND sg13g2_decap_8
X_4529_ VGND VPWR _1479_ _1478_ _1477_ sg13g2_or2_1
Xhold230 _0232_ VPWR VGND net882 sg13g2_dlygate4sd3_1
XFILLER_49_14 VPWR VGND sg13g2_decap_8
Xhold263 ppwm_i.u_ppwm.u_mem.memory\[52\] VPWR VGND net915 sg13g2_dlygate4sd3_1
XFILLER_46_1028 VPWR VGND sg13g2_fill_1
Xhold296 ppwm_i.u_ppwm.u_mem.memory\[81\] VPWR VGND net948 sg13g2_dlygate4sd3_1
Xhold285 falu_i.falutop.div_inst.val\[5\] VPWR VGND net937 sg13g2_dlygate4sd3_1
Xhold274 falu_i.falutop.i2c_inst.data_in\[12\] VPWR VGND net926 sg13g2_dlygate4sd3_1
Xfanout721 net722 net721 VPWR VGND sg13g2_buf_8
Xfanout710 net715 net710 VPWR VGND sg13g2_buf_8
Xfanout732 net733 net732 VPWR VGND sg13g2_buf_8
Xfanout743 net746 net743 VPWR VGND sg13g2_buf_8
Xfanout776 net1178 net776 VPWR VGND sg13g2_buf_8
Xfanout754 falu_i.falutop.alu_data_in\[4\] net754 VPWR VGND sg13g2_buf_8
Xfanout765 falu_i.falutop.alu_data_in\[2\] net765 VPWR VGND sg13g2_buf_8
XFILLER_46_616 VPWR VGND sg13g2_decap_8
Xfanout787 ppwm_i.u_ppwm.pc\[3\] net787 VPWR VGND sg13g2_buf_1
Xfanout798 net799 net798 VPWR VGND sg13g2_buf_8
XFILLER_42_800 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_41_376 VPWR VGND sg13g2_decap_8
XFILLER_14_579 VPWR VGND sg13g2_fill_2
XFILLER_6_723 VPWR VGND sg13g2_decap_8
XFILLER_6_778 VPWR VGND sg13g2_fill_2
XFILLER_7_1000 VPWR VGND sg13g2_decap_8
XFILLER_2_995 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_4
X_5499__277 VPWR VGND net277 sg13g2_tiehi
XFILLER_18_830 VPWR VGND sg13g2_decap_8
XFILLER_36_126 VPWR VGND sg13g2_fill_1
X_3900_ VGND VPWR _2186_ net670 _0169_ _0978_ sg13g2_a21oi_1
X_4880_ _1825_ _1790_ _1823_ VPWR VGND sg13g2_xnor2_1
X_3831_ net829 VPWR _0944_ VGND ppwm_i.u_ppwm.u_mem.memory\[36\] net643 sg13g2_o21ai_1
XFILLER_32_354 VPWR VGND sg13g2_fill_2
X_3762_ VGND VPWR _2234_ net662 _0100_ _0909_ sg13g2_a21oi_1
X_5501_ net273 VGND VPWR _0260_ falu_i.falutop.div_inst.b1\[5\] clknet_leaf_2_clk
+ sg13g2_dfrbpq_1
X_3693_ _0722_ net569 _0854_ _0855_ VPWR VGND sg13g2_nor3_1
X_5432_ net163 VGND VPWR net391 ppwm_i.u_ppwm.u_mem.memory\[91\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_5363_ net326 VGND VPWR _0122_ ppwm_i.u_ppwm.u_mem.memory\[22\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_4314_ VGND VPWR _1235_ _1266_ _1267_ _1265_ sg13g2_a21oi_1
X_5294_ net109 VGND VPWR net956 ppwm_i.u_ppwm.global_counter\[11\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_4245_ _1206_ net498 net607 VPWR VGND sg13g2_nand2_1
X_4176_ net819 VPWR _1153_ VGND falu_i.falutop.div_inst.val\[7\] net637 sg13g2_o21ai_1
X_3127_ VGND VPWR net802 _0361_ _0012_ _0362_ sg13g2_a21oi_1
XFILLER_27_148 VPWR VGND sg13g2_fill_1
X_5374__304 VPWR VGND net304 sg13g2_tiehi
X_3058_ _2412_ _2203_ net692 VPWR VGND sg13g2_nand2_1
XFILLER_36_660 VPWR VGND sg13g2_decap_8
XFILLER_36_682 VPWR VGND sg13g2_fill_1
XFILLER_23_310 VPWR VGND sg13g2_fill_2
XFILLER_24_844 VPWR VGND sg13g2_decap_8
XFILLER_13_1027 VPWR VGND sg13g2_fill_2
XFILLER_3_737 VPWR VGND sg13g2_fill_1
Xfanout573 _0615_ net573 VPWR VGND sg13g2_buf_8
Xfanout584 net585 net584 VPWR VGND sg13g2_buf_8
XFILLER_47_925 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_4
Xfanout595 net596 net595 VPWR VGND sg13g2_buf_1
XFILLER_46_457 VPWR VGND sg13g2_fill_1
XFILLER_46_446 VPWR VGND sg13g2_decap_8
XFILLER_34_608 VPWR VGND sg13g2_decap_8
XFILLER_15_800 VPWR VGND sg13g2_fill_1
XFILLER_15_833 VPWR VGND sg13g2_decap_8
XFILLER_14_398 VPWR VGND sg13g2_decap_4
XFILLER_10_571 VPWR VGND sg13g2_fill_1
XFILLER_6_542 VPWR VGND sg13g2_decap_4
XFILLER_10_593 VPWR VGND sg13g2_decap_8
XFILLER_29_1012 VPWR VGND sg13g2_decap_8
XFILLER_49_251 VPWR VGND sg13g2_decap_8
XFILLER_2_20 VPWR VGND sg13g2_fill_1
X_4030_ net1043 _1049_ _1056_ VPWR VGND sg13g2_nor2_1
XFILLER_2_86 VPWR VGND sg13g2_fill_1
XFILLER_18_671 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_44_clk clknet_3_0__leaf_clk clknet_leaf_44_clk VPWR VGND sg13g2_buf_8
X_4932_ _1876_ _1842_ _1875_ VPWR VGND sg13g2_xnor2_1
XFILLER_24_129 VPWR VGND sg13g2_decap_8
X_4863_ _1761_ VPWR _1808_ VGND _1759_ _1762_ sg13g2_o21ai_1
XFILLER_20_324 VPWR VGND sg13g2_decap_8
XFILLER_21_847 VPWR VGND sg13g2_decap_8
XFILLER_32_162 VPWR VGND sg13g2_fill_2
X_4794_ _1704_ VPWR _1740_ VGND _1685_ _1705_ sg13g2_o21ai_1
XFILLER_20_357 VPWR VGND sg13g2_fill_2
X_3814_ VGND VPWR _2216_ net641 _0126_ _0935_ sg13g2_a21oi_1
X_3745_ _0901_ net459 net1015 VPWR VGND sg13g2_nand2_1
XFILLER_21_29 VPWR VGND sg13g2_fill_2
X_5415_ net222 VGND VPWR net384 ppwm_i.u_ppwm.u_mem.memory\[74\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_3676_ _2240_ net586 _0839_ VPWR VGND sg13g2_nor2_1
X_5346_ net360 VGND VPWR net484 ppwm_i.u_ppwm.u_mem.memory\[5\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_5277_ net142 VGND VPWR net1061 ppwm_i.u_ppwm.u_pwm.counter\[5\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_2
X_4228_ VGND VPWR net605 _1192_ _0282_ _1193_ sg13g2_a21oi_1
X_4159_ falu_i.falutop.div_inst.b1\[7\] net1054 _1103_ _0262_ VPWR VGND sg13g2_mux2_1
XFILLER_15_107 VPWR VGND sg13g2_fill_2
XFILLER_43_438 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_35_clk clknet_3_5__leaf_clk clknet_leaf_35_clk VPWR VGND sg13g2_buf_8
XFILLER_23_173 VPWR VGND sg13g2_fill_1
XFILLER_3_578 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_fill_1
XFILLER_46_254 VPWR VGND sg13g2_decap_8
XFILLER_28_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_26_clk clknet_3_6__leaf_clk clknet_leaf_26_clk VPWR VGND sg13g2_buf_8
XFILLER_43_961 VPWR VGND sg13g2_decap_8
XFILLER_15_674 VPWR VGND sg13g2_fill_1
X_5468__349 VPWR VGND net349 sg13g2_tiehi
X_3530_ _0703_ ppwm_i.u_ppwm.global_counter\[13\] net593 VPWR VGND sg13g2_nand2_1
XFILLER_7_895 VPWR VGND sg13g2_decap_8
X_5583__231 VPWR VGND net231 sg13g2_tiehi
X_3461_ VGND VPWR _0637_ _0616_ net579 sg13g2_or2_1
X_3392_ VPWR VGND _0569_ net610 _0566_ _0547_ _0570_ _0549_ sg13g2_a221oi_1
X_5200_ net967 net623 _2116_ VPWR VGND sg13g2_nor2_1
X_5131_ _1834_ VPWR _2070_ VGND _2068_ _2069_ sg13g2_o21ai_1
X_5062_ _2003_ _2002_ _2001_ VPWR VGND sg13g2_nand2b_1
X_4013_ ppwm_i.u_ppwm.u_mem.bit_count\[5\] net806 _1043_ VPWR VGND net512 sg13g2_nand3b_1
XFILLER_16_18 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_17_clk clknet_3_4__leaf_clk clknet_leaf_17_clk VPWR VGND sg13g2_buf_8
Xheichips25_tiny_wrapper_9 VPWR VGND uio_oe[1] sg13g2_tielo
X_4915_ net719 net712 net761 net758 _1859_ VPWR VGND sg13g2_and4_1
XFILLER_34_983 VPWR VGND sg13g2_decap_8
X_4846_ VGND VPWR _1742_ _1745_ _1791_ _1743_ sg13g2_a21oi_1
X_4777_ _1722_ VPWR _1723_ VGND _1660_ _1663_ sg13g2_o21ai_1
X_3728_ net602 net783 _0886_ VPWR VGND sg13g2_xor2_1
X_3659_ VGND VPWR _0824_ _0823_ _0815_ sg13g2_or2_1
XFILLER_0_504 VPWR VGND sg13g2_decap_8
X_5329_ net43 VGND VPWR _0088_ ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] clknet_leaf_17_clk
+ sg13g2_dfrbpq_2
XFILLER_0_548 VPWR VGND sg13g2_fill_1
XFILLER_28_210 VPWR VGND sg13g2_decap_8
XFILLER_28_232 VPWR VGND sg13g2_fill_2
XFILLER_16_405 VPWR VGND sg13g2_decap_4
XFILLER_17_939 VPWR VGND sg13g2_decap_8
XFILLER_28_298 VPWR VGND sg13g2_decap_4
XFILLER_40_953 VPWR VGND sg13g2_decap_8
XFILLER_12_633 VPWR VGND sg13g2_fill_1
XFILLER_4_887 VPWR VGND sg13g2_decap_8
X_5400__252 VPWR VGND net252 sg13g2_tiehi
XFILLER_34_257 VPWR VGND sg13g2_fill_1
XFILLER_16_972 VPWR VGND sg13g2_decap_8
X_2961_ VPWR VGND _2165_ net708 net694 _2174_ _2315_ net697 sg13g2_a221oi_1
X_4700_ VPWR VGND _1647_ _1075_ _1646_ net614 _1648_ _1643_ sg13g2_a221oi_1
X_2892_ net1187 _2246_ VPWR VGND sg13g2_inv_4
X_4631_ _1263_ _1269_ _1239_ _1580_ VPWR VGND sg13g2_nand3_1
XFILLER_30_463 VPWR VGND sg13g2_fill_2
XFILLER_31_975 VPWR VGND sg13g2_decap_8
X_4562_ VPWR VGND _1510_ _1511_ _1509_ _1225_ _1512_ _1383_ sg13g2_a221oi_1
X_4493_ _1444_ _1230_ _1427_ VPWR VGND sg13g2_xnor2_1
X_3513_ _0686_ VPWR _0687_ VGND net1171 _0614_ sg13g2_o21ai_1
X_3444_ _0620_ _0616_ _2344_ VPWR VGND sg13g2_nand2b_1
Xclkbuf_leaf_6_clk clknet_3_1__leaf_clk clknet_leaf_6_clk VPWR VGND sg13g2_buf_8
XFILLER_40_0 VPWR VGND sg13g2_decap_8
X_3375_ _0553_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] ppwm_i.u_ppwm.global_counter\[0\]
+ VPWR VGND sg13g2_nand2b_1
X_5114_ VGND VPWR _2009_ _2039_ _2053_ _2052_ sg13g2_a21oi_1
X_5045_ _1956_ _1958_ _1986_ VPWR VGND sg13g2_nor2_1
Xheichips25_tiny_wrapper_12 VPWR VGND uio_oe[4] sg13g2_tielo
Xheichips25_tiny_wrapper_23 VPWR VGND uio_out[7] sg13g2_tielo
X_5260__175 VPWR VGND net175 sg13g2_tiehi
XFILLER_25_213 VPWR VGND sg13g2_decap_4
XFILLER_25_246 VPWR VGND sg13g2_fill_1
XFILLER_22_964 VPWR VGND sg13g2_decap_8
X_4829_ _1775_ _1740_ _1773_ VPWR VGND sg13g2_xnor2_1
XFILLER_0_312 VPWR VGND sg13g2_fill_1
X_5382__288 VPWR VGND net288 sg13g2_tiehi
XFILLER_1_868 VPWR VGND sg13g2_decap_8
XFILLER_49_839 VPWR VGND sg13g2_fill_2
XFILLER_16_202 VPWR VGND sg13g2_fill_2
XFILLER_17_747 VPWR VGND sg13g2_fill_1
XFILLER_16_235 VPWR VGND sg13g2_fill_1
XFILLER_17_61 VPWR VGND sg13g2_fill_2
XFILLER_17_72 VPWR VGND sg13g2_fill_2
XFILLER_9_902 VPWR VGND sg13g2_decap_8
XFILLER_12_463 VPWR VGND sg13g2_fill_1
XFILLER_13_964 VPWR VGND sg13g2_decap_8
XFILLER_9_979 VPWR VGND sg13g2_decap_8
X_5283__131 VPWR VGND net131 sg13g2_tiehi
XFILLER_39_316 VPWR VGND sg13g2_decap_8
X_3160_ ppwm_i.u_ppwm.u_pwm.counter\[3\] ppwm_i.u_ppwm.u_pwm.counter\[2\] ppwm_i.u_ppwm.u_pwm.counter\[1\]
+ ppwm_i.u_ppwm.u_pwm.counter\[0\] _0384_ VPWR VGND sg13g2_nor4_1
XFILLER_39_349 VPWR VGND sg13g2_fill_2
XFILLER_39_327 VPWR VGND sg13g2_fill_2
XFILLER_0_890 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_8
X_3091_ net985 _2440_ _2441_ VPWR VGND sg13g2_nor2b_1
Xhold1 ppwm_i.u_ppwm.u_mem.data_sync1 VPWR VGND net373 sg13g2_dlygate4sd3_1
XFILLER_48_872 VPWR VGND sg13g2_decap_8
XFILLER_23_706 VPWR VGND sg13g2_decap_8
X_3993_ net808 _1027_ _0213_ VPWR VGND sg13g2_and2_1
X_2944_ VPWR _2298_ net877 VGND sg13g2_inv_1
X_2875_ VPWR _2229_ net441 VGND sg13g2_inv_1
X_4614_ _1563_ _1548_ _1562_ VPWR VGND sg13g2_nand2b_1
X_4545_ _1495_ _1431_ _1493_ VPWR VGND sg13g2_xnor2_1
Xhold401 _0214_ VPWR VGND net1053 sg13g2_dlygate4sd3_1
Xhold434 falu_i.falutop.data_in\[13\] VPWR VGND net1086 sg13g2_dlygate4sd3_1
Xhold412 falu_i.falutop.i2c_inst.result\[9\] VPWR VGND net1064 sg13g2_dlygate4sd3_1
Xhold423 _2101_ VPWR VGND net1075 sg13g2_dlygate4sd3_1
Xhold445 falu_i.falutop.i2c_inst.counter\[2\] VPWR VGND net1097 sg13g2_dlygate4sd3_1
Xhold467 falu_i.falutop.div_inst.rem\[3\] VPWR VGND net1119 sg13g2_dlygate4sd3_1
X_4476_ VGND VPWR _1219_ _1234_ _1427_ _1232_ sg13g2_a21oi_1
Xhold478 _0447_ VPWR VGND net1130 sg13g2_dlygate4sd3_1
Xhold456 _0432_ VPWR VGND net1108 sg13g2_dlygate4sd3_1
X_3427_ _0604_ net1162 _0516_ _0605_ VPWR VGND sg13g2_mux2_1
Xhold489 falu_i.falutop.data_in\[1\] VPWR VGND net1141 sg13g2_dlygate4sd3_1
X_3358_ _0536_ net784 ppwm_i.u_ppwm.global_counter\[1\] VPWR VGND sg13g2_nand2b_1
X_3289_ VGND VPWR _2274_ ppwm_i.u_ppwm.u_pwm.cmp_value\[8\] _0472_ _0471_ sg13g2_a21oi_1
X_5028_ _1969_ VPWR _1970_ VGND net731 net563 sg13g2_o21ai_1
XFILLER_14_717 VPWR VGND sg13g2_decap_4
XFILLER_10_901 VPWR VGND sg13g2_decap_8
XFILLER_16_1014 VPWR VGND sg13g2_decap_8
XFILLER_6_927 VPWR VGND sg13g2_decap_8
XFILLER_10_978 VPWR VGND sg13g2_decap_8
XFILLER_49_625 VPWR VGND sg13g2_decap_8
XFILLER_1_698 VPWR VGND sg13g2_fill_2
XFILLER_37_809 VPWR VGND sg13g2_fill_2
XFILLER_36_319 VPWR VGND sg13g2_decap_8
XFILLER_17_599 VPWR VGND sg13g2_decap_8
XFILLER_13_794 VPWR VGND sg13g2_decap_8
XFILLER_5_993 VPWR VGND sg13g2_decap_8
X_4330_ net770 net744 net566 _1283_ VPWR VGND sg13g2_mux2_1
X_4261_ _2296_ _2305_ _1214_ VPWR VGND sg13g2_nor2_2
X_3212_ ppwm_i.u_ppwm.u_pwm.counter\[7\] _0415_ net1094 _0418_ VPWR VGND sg13g2_nand3_1
X_4192_ _1165_ _1121_ _1122_ VPWR VGND sg13g2_xnor2_1
X_5320__61 VPWR VGND net61 sg13g2_tiehi
X_3143_ VGND VPWR net802 _0372_ _0017_ _0373_ sg13g2_a21oi_1
X_3074_ net386 VPWR _0001_ VGND _2421_ _2422_ sg13g2_o21ai_1
XFILLER_36_831 VPWR VGND sg13g2_fill_2
XFILLER_35_352 VPWR VGND sg13g2_fill_2
XFILLER_23_547 VPWR VGND sg13g2_fill_2
XFILLER_23_569 VPWR VGND sg13g2_decap_8
X_3976_ VGND VPWR _2159_ net648 _0207_ _1016_ sg13g2_a21oi_1
X_2927_ _2281_ net430 VPWR VGND sg13g2_inv_2
XFILLER_10_208 VPWR VGND sg13g2_fill_1
XFILLER_31_591 VPWR VGND sg13g2_decap_8
X_2858_ VPWR _2212_ net534 VGND sg13g2_inv_1
X_5577_ net307 VGND VPWR net907 falu_i.falutop.div_inst.a\[0\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_1
Xhold220 _0235_ VPWR VGND net872 sg13g2_dlygate4sd3_1
Xhold253 falu_i.falutop.div_inst.val\[4\] VPWR VGND net905 sg13g2_dlygate4sd3_1
X_4528_ _1478_ _1423_ _1425_ VPWR VGND sg13g2_nand2_1
Xhold242 falu_i.falutop.i2c_inst.data_in\[13\] VPWR VGND net894 sg13g2_dlygate4sd3_1
Xhold231 ppwm_i.u_ppwm.u_mem.programming VPWR VGND net883 sg13g2_dlygate4sd3_1
XFILLER_46_1007 VPWR VGND sg13g2_decap_8
Xhold264 _0151_ VPWR VGND net916 sg13g2_dlygate4sd3_1
X_4459_ VPWR _1410_ _1409_ VGND sg13g2_inv_1
Xhold275 _0240_ VPWR VGND net927 sg13g2_dlygate4sd3_1
Xhold286 falu_i.falutop.alu_inst.op\[2\] VPWR VGND net938 sg13g2_dlygate4sd3_1
Xfanout700 net701 net700 VPWR VGND sg13g2_buf_8
Xhold297 ppwm_i.u_ppwm.u_mem.memory\[47\] VPWR VGND net949 sg13g2_dlygate4sd3_1
Xfanout711 net713 net711 VPWR VGND sg13g2_buf_8
Xfanout722 falu_i.falutop.alu_data_in\[13\] net722 VPWR VGND sg13g2_buf_2
Xfanout733 net734 net733 VPWR VGND sg13g2_buf_8
Xfanout755 net758 net755 VPWR VGND sg13g2_buf_2
Xfanout744 net746 net744 VPWR VGND sg13g2_buf_8
Xfanout766 net767 net766 VPWR VGND sg13g2_buf_8
Xfanout788 net790 net788 VPWR VGND sg13g2_buf_8
Xfanout777 falu_i.falutop.data_in\[7\] net777 VPWR VGND sg13g2_buf_8
Xfanout799 _2294_ net799 VPWR VGND sg13g2_buf_8
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_41_300 VPWR VGND sg13g2_decap_4
XFILLER_10_797 VPWR VGND sg13g2_decap_8
XFILLER_5_234 VPWR VGND sg13g2_decap_4
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_2_974 VPWR VGND sg13g2_decap_8
XFILLER_1_451 VPWR VGND sg13g2_fill_2
XFILLER_49_455 VPWR VGND sg13g2_decap_8
X_5448__98 VPWR VGND net98 sg13g2_tiehi
XFILLER_18_886 VPWR VGND sg13g2_decap_8
X_3830_ VGND VPWR _2210_ net656 _0134_ _0943_ sg13g2_a21oi_1
X_3761_ net836 VPWR _0909_ VGND net868 net662 sg13g2_o21ai_1
XFILLER_9_540 VPWR VGND sg13g2_fill_1
X_5500_ net275 VGND VPWR _0259_ falu_i.falutop.div_inst.b1\[4\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_3692_ VGND VPWR net581 _0724_ _0854_ _0853_ sg13g2_a21oi_1
X_5431_ net167 VGND VPWR net958 ppwm_i.u_ppwm.u_mem.memory\[90\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_5362_ net328 VGND VPWR net478 ppwm_i.u_ppwm.u_mem.memory\[21\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_4313_ _1266_ net745 _2301_ VPWR VGND sg13g2_nand2_1
X_5293_ net111 VGND VPWR _0055_ ppwm_i.u_ppwm.global_counter\[10\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_4244_ VGND VPWR net606 _1204_ _0286_ _1205_ sg13g2_a21oi_1
X_4175_ VGND VPWR _2147_ net637 _0270_ _1152_ sg13g2_a21oi_1
X_5478__329 VPWR VGND net329 sg13g2_tiehi
XFILLER_28_606 VPWR VGND sg13g2_fill_1
X_3126_ net804 VPWR _0362_ VGND net873 _0361_ sg13g2_o21ai_1
X_3057_ VGND VPWR _2208_ net688 _2411_ net708 sg13g2_a21oi_1
XFILLER_24_823 VPWR VGND sg13g2_decap_8
XFILLER_13_1006 VPWR VGND sg13g2_decap_8
X_3959_ net837 VPWR _1008_ VGND ppwm_i.u_ppwm.u_mem.memory\[100\] net648 sg13g2_o21ai_1
XFILLER_3_727 VPWR VGND sg13g2_fill_2
XFILLER_3_705 VPWR VGND sg13g2_decap_8
XFILLER_3_749 VPWR VGND sg13g2_decap_8
XFILLER_2_215 VPWR VGND sg13g2_fill_1
XFILLER_2_248 VPWR VGND sg13g2_fill_1
XFILLER_47_904 VPWR VGND sg13g2_decap_8
Xfanout574 _0649_ net574 VPWR VGND sg13g2_buf_8
Xfanout563 net564 net563 VPWR VGND sg13g2_buf_8
Xfanout585 _2390_ net585 VPWR VGND sg13g2_buf_1
Xfanout596 net597 net596 VPWR VGND sg13g2_buf_8
XFILLER_42_664 VPWR VGND sg13g2_fill_1
XFILLER_15_889 VPWR VGND sg13g2_decap_8
XFILLER_25_72 VPWR VGND sg13g2_fill_1
XFILLER_30_837 VPWR VGND sg13g2_fill_2
XFILLER_10_583 VPWR VGND sg13g2_decap_4
XFILLER_49_230 VPWR VGND sg13g2_decap_8
XFILLER_2_76 VPWR VGND sg13g2_fill_1
XFILLER_45_480 VPWR VGND sg13g2_fill_2
X_4931_ _1875_ _1872_ _1874_ VPWR VGND sg13g2_nand2_1
XFILLER_17_171 VPWR VGND sg13g2_decap_8
X_4862_ _1806_ _1801_ _1807_ VPWR VGND sg13g2_xor2_1
XFILLER_33_642 VPWR VGND sg13g2_fill_2
XFILLER_21_826 VPWR VGND sg13g2_decap_8
XFILLER_32_152 VPWR VGND sg13g2_fill_1
XFILLER_32_174 VPWR VGND sg13g2_fill_1
X_3813_ net824 VPWR _0935_ VGND net963 net641 sg13g2_o21ai_1
XFILLER_33_697 VPWR VGND sg13g2_decap_8
X_4793_ VGND VPWR _1679_ _1711_ _1739_ _1710_ sg13g2_a21oi_1
X_3744_ VPWR VGND _0900_ net798 _0897_ _2235_ _0091_ net570 sg13g2_a221oi_1
X_5410__232 VPWR VGND net232 sg13g2_tiehi
X_3675_ _0832_ VPWR _0838_ VGND _2241_ net586 sg13g2_o21ai_1
X_5414_ net224 VGND VPWR net923 ppwm_i.u_ppwm.u_mem.memory\[73\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_5345_ net362 VGND VPWR _0104_ ppwm_i.u_ppwm.u_mem.memory\[4\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_5276_ net144 VGND VPWR net1091 ppwm_i.u_ppwm.u_pwm.counter\[4\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_2
X_4227_ net435 net605 _1193_ VPWR VGND sg13g2_nor2_1
XFILLER_46_38 VPWR VGND sg13g2_fill_2
X_4158_ net1056 net920 _1103_ _0261_ VPWR VGND sg13g2_mux2_1
XFILLER_43_406 VPWR VGND sg13g2_fill_1
X_5558__194 VPWR VGND net194 sg13g2_tiehi
XFILLER_16_609 VPWR VGND sg13g2_decap_4
X_3109_ net985 _2154_ _0349_ VPWR VGND sg13g2_nor2_1
X_4089_ VPWR VGND net986 _1092_ _1091_ net985 _1093_ _1084_ sg13g2_a221oi_1
XFILLER_37_992 VPWR VGND sg13g2_decap_8
XFILLER_24_631 VPWR VGND sg13g2_decap_8
XFILLER_24_664 VPWR VGND sg13g2_decap_8
XFILLER_24_697 VPWR VGND sg13g2_decap_8
XFILLER_20_881 VPWR VGND sg13g2_decap_8
XFILLER_46_200 VPWR VGND sg13g2_fill_2
X_5392__268 VPWR VGND net268 sg13g2_tiehi
XFILLER_43_940 VPWR VGND sg13g2_decap_8
XFILLER_36_93 VPWR VGND sg13g2_fill_1
XFILLER_14_174 VPWR VGND sg13g2_decap_4
XFILLER_30_689 VPWR VGND sg13g2_fill_2
XFILLER_11_881 VPWR VGND sg13g2_decap_8
XFILLER_7_874 VPWR VGND sg13g2_decap_8
XFILLER_6_373 VPWR VGND sg13g2_fill_2
X_3460_ _0636_ net571 _0635_ _0627_ _0622_ VPWR VGND sg13g2_a22oi_1
X_3391_ _0565_ _0568_ _0569_ VPWR VGND sg13g2_nor2_1
X_5130_ _1281_ VPWR _2069_ VGND net717 net563 sg13g2_o21ai_1
X_5061_ _2002_ _1986_ _2000_ VPWR VGND sg13g2_nand2_1
X_4012_ _1042_ net512 _1040_ VPWR VGND sg13g2_nand2_1
XFILLER_38_789 VPWR VGND sg13g2_fill_1
XFILLER_38_767 VPWR VGND sg13g2_fill_1
XFILLER_37_255 VPWR VGND sg13g2_fill_2
X_5293__111 VPWR VGND net111 sg13g2_tiehi
X_4914_ _1858_ net758 net718 net761 net712 VPWR VGND sg13g2_a22oi_1
XFILLER_34_962 VPWR VGND sg13g2_decap_8
X_4845_ _1770_ VPWR _1790_ VGND _1748_ _1771_ sg13g2_o21ai_1
XFILLER_32_18 VPWR VGND sg13g2_fill_2
X_4776_ _1722_ _1719_ _1720_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_133 VPWR VGND sg13g2_fill_2
X_3727_ _0885_ net783 net602 VPWR VGND sg13g2_nand2_1
X_3658_ _0823_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] net611 VPWR VGND sg13g2_xnor2_1
X_3589_ _0759_ _0756_ _0758_ VPWR VGND sg13g2_nand2_1
X_5328_ net45 VGND VPWR net1175 ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
XFILLER_0_527 VPWR VGND sg13g2_fill_1
X_5259_ net177 VGND VPWR _0021_ falu_i.falutop.i2c_inst.data_in\[17\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
XFILLER_44_715 VPWR VGND sg13g2_fill_2
XFILLER_17_918 VPWR VGND sg13g2_decap_8
XFILLER_43_225 VPWR VGND sg13g2_decap_8
XFILLER_43_236 VPWR VGND sg13g2_fill_2
XFILLER_25_995 VPWR VGND sg13g2_decap_8
XFILLER_40_932 VPWR VGND sg13g2_decap_8
XFILLER_11_111 VPWR VGND sg13g2_fill_1
XFILLER_4_866 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_39_509 VPWR VGND sg13g2_decap_8
XFILLER_19_200 VPWR VGND sg13g2_fill_1
XFILLER_16_951 VPWR VGND sg13g2_decap_8
X_2960_ _2314_ net690 _2170_ net702 _2160_ VPWR VGND sg13g2_a22oi_1
X_2891_ _2245_ net1190 VPWR VGND sg13g2_inv_2
XFILLER_31_954 VPWR VGND sg13g2_decap_8
X_4630_ _1500_ _1573_ _1578_ _1579_ VPWR VGND sg13g2_nor3_1
XFILLER_33_1009 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_fill_1
X_4561_ _1225_ _1323_ _1511_ VPWR VGND sg13g2_nor2_1
X_4492_ _1442_ VPWR _1443_ VGND _1228_ _1319_ sg13g2_o21ai_1
X_3512_ _0679_ _0685_ _0672_ _0686_ VPWR VGND sg13g2_nand3_1
X_3443_ _0619_ ppwm_i.u_ppwm.pwm_value\[0\] net608 VPWR VGND sg13g2_nand2_1
X_5113_ _2042_ VPWR _2052_ VGND _2037_ _2038_ sg13g2_o21ai_1
X_3374_ _0552_ _2240_ ppwm_i.u_ppwm.global_counter\[3\] VPWR VGND sg13g2_nand2_1
X_5044_ _1941_ VPWR _1985_ VGND _1897_ _1942_ sg13g2_o21ai_1
Xheichips25_tiny_wrapper_13 VPWR VGND uio_oe[5] sg13g2_tielo
XFILLER_38_553 VPWR VGND sg13g2_fill_1
XFILLER_38_542 VPWR VGND sg13g2_fill_2
Xheichips25_tiny_wrapper_24 VPWR VGND uo_out[1] sg13g2_tielo
XFILLER_38_597 VPWR VGND sg13g2_fill_1
XFILLER_22_943 VPWR VGND sg13g2_decap_8
X_4828_ _1774_ _1740_ _1773_ VPWR VGND sg13g2_nand2_1
XFILLER_21_464 VPWR VGND sg13g2_decap_4
XFILLER_5_619 VPWR VGND sg13g2_fill_2
X_4759_ _1703_ _1686_ _1706_ VPWR VGND sg13g2_xor2_1
XFILLER_49_1027 VPWR VGND sg13g2_fill_2
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_17_715 VPWR VGND sg13g2_decap_4
XFILLER_13_943 VPWR VGND sg13g2_decap_8
XFILLER_9_958 VPWR VGND sg13g2_decap_8
X_5572__48 VPWR VGND net48 sg13g2_tiehi
XFILLER_4_641 VPWR VGND sg13g2_decap_8
X_5545__355 VPWR VGND net355 sg13g2_tiehi
X_3090_ net1097 falu_i.falutop.i2c_inst.counter\[1\] net1045 _2440_ VPWR VGND sg13g2_nor3_1
Xhold2 ppwm_i.u_ppwm.u_mem.clk_prog_sync1 VPWR VGND net374 sg13g2_dlygate4sd3_1
XFILLER_48_851 VPWR VGND sg13g2_decap_8
XFILLER_47_383 VPWR VGND sg13g2_fill_1
X_3992_ _1024_ VPWR _1027_ VGND _1025_ _1026_ sg13g2_o21ai_1
X_2943_ net716 _2297_ VPWR VGND sg13g2_inv_4
X_2874_ VPWR _2228_ net504 VGND sg13g2_inv_1
X_4613_ _1562_ _1552_ _1561_ VPWR VGND sg13g2_xnor2_1
Xhold402 falu_i.falutop.div_inst.b\[7\] VPWR VGND net1054 sg13g2_dlygate4sd3_1
X_4544_ VGND VPWR _1494_ _1493_ _1432_ sg13g2_or2_1
Xhold424 ppwm_i.u_ppwm.global_counter\[18\] VPWR VGND net1076 sg13g2_dlygate4sd3_1
Xhold435 _0326_ VPWR VGND net1087 sg13g2_dlygate4sd3_1
Xhold413 _0304_ VPWR VGND net1065 sg13g2_dlygate4sd3_1
X_4475_ VGND VPWR _1399_ _1424_ _1426_ _1310_ sg13g2_a21oi_1
Xhold446 falu_i.falutop.div_inst.rem\[1\] VPWR VGND net1098 sg13g2_dlygate4sd3_1
Xhold468 ppwm_i.u_ppwm.global_counter\[10\] VPWR VGND net1120 sg13g2_dlygate4sd3_1
Xhold457 _0049_ VPWR VGND net1109 sg13g2_dlygate4sd3_1
X_3426_ _0532_ VPWR _0604_ VGND _0570_ _0603_ sg13g2_o21ai_1
Xhold479 falu_i.falutop.alu_data_in\[6\] VPWR VGND net1131 sg13g2_dlygate4sd3_1
X_3357_ _0534_ ppwm_i.u_ppwm.pwm_value\[0\] _0535_ VPWR VGND ppwm_i.u_ppwm.global_counter\[0\]
+ sg13g2_nand3b_1
XFILLER_38_17 VPWR VGND sg13g2_decap_8
X_3288_ _0470_ VPWR _0471_ VGND ppwm_i.u_ppwm.u_pwm.counter\[7\] _2281_ sg13g2_o21ai_1
XFILLER_39_840 VPWR VGND sg13g2_decap_8
X_5027_ _1969_ net563 net760 VPWR VGND sg13g2_nand2b_1
XFILLER_14_729 VPWR VGND sg13g2_fill_2
XFILLER_22_740 VPWR VGND sg13g2_fill_1
XFILLER_6_906 VPWR VGND sg13g2_decap_8
XFILLER_10_957 VPWR VGND sg13g2_decap_8
XFILLER_1_633 VPWR VGND sg13g2_fill_2
XFILLER_49_604 VPWR VGND sg13g2_fill_1
XFILLER_48_125 VPWR VGND sg13g2_fill_2
XFILLER_49_659 VPWR VGND sg13g2_fill_1
X_5575__359 VPWR VGND net359 sg13g2_tiehi
XFILLER_28_83 VPWR VGND sg13g2_fill_1
XFILLER_45_865 VPWR VGND sg13g2_fill_2
XFILLER_17_523 VPWR VGND sg13g2_decap_4
XFILLER_44_375 VPWR VGND sg13g2_fill_1
XFILLER_12_250 VPWR VGND sg13g2_fill_2
XFILLER_9_766 VPWR VGND sg13g2_fill_1
XFILLER_5_972 VPWR VGND sg13g2_decap_8
X_4260_ VPWR _0294_ net880 VGND sg13g2_inv_1
XFILLER_5_98 VPWR VGND sg13g2_decap_4
X_3211_ _0041_ net809 _0416_ _0417_ VPWR VGND sg13g2_and3_1
X_4191_ VGND VPWR net633 _1163_ _0274_ _1164_ sg13g2_a21oi_1
X_3142_ net816 VPWR _0373_ VGND net894 _0372_ sg13g2_o21ai_1
XFILLER_39_136 VPWR VGND sg13g2_decap_8
X_3073_ net821 net385 _2426_ VPWR VGND ppwm_i.u_ppwm.period_start sg13g2_nand3b_1
XFILLER_48_692 VPWR VGND sg13g2_fill_1
XFILLER_36_843 VPWR VGND sg13g2_fill_2
XFILLER_39_1015 VPWR VGND sg13g2_decap_8
X_3975_ net838 VPWR _1016_ VGND net540 net648 sg13g2_o21ai_1
X_2926_ VPWR _2280_ net924 VGND sg13g2_inv_1
X_2857_ VPWR _2211_ net547 VGND sg13g2_inv_1
Xhold210 _0242_ VPWR VGND net862 sg13g2_dlygate4sd3_1
X_5576_ net351 VGND VPWR net921 falu_i.falutop.div_inst.b\[6\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4527_ _1476_ _1462_ _1477_ VPWR VGND sg13g2_xor2_1
Xhold243 _0241_ VPWR VGND net895 sg13g2_dlygate4sd3_1
Xhold221 falu_i.falutop.i2c_inst.data_in\[8\] VPWR VGND net873 sg13g2_dlygate4sd3_1
Xhold232 _0907_ VPWR VGND net884 sg13g2_dlygate4sd3_1
Xhold287 falu_i.falutop.div_inst.val\[1\] VPWR VGND net939 sg13g2_dlygate4sd3_1
Xhold254 falu_i.falutop.div_inst.a\[0\] VPWR VGND net906 sg13g2_dlygate4sd3_1
Xhold265 falu_i.falutop.div_inst.i\[1\] VPWR VGND net917 sg13g2_dlygate4sd3_1
X_4458_ VGND VPWR _1409_ _1358_ _1353_ sg13g2_or2_1
Xhold276 ppwm_i.u_ppwm.u_mem.memory\[14\] VPWR VGND net928 sg13g2_dlygate4sd3_1
X_3409_ _0587_ _2235_ ppwm_i.u_ppwm.global_counter\[19\] VPWR VGND sg13g2_nand2_1
Xfanout723 net724 net723 VPWR VGND sg13g2_buf_8
Xfanout712 net713 net712 VPWR VGND sg13g2_buf_1
Xhold298 ppwm_i.u_ppwm.u_mem.memory\[25\] VPWR VGND net950 sg13g2_dlygate4sd3_1
Xfanout701 net704 net701 VPWR VGND sg13g2_buf_8
X_4389_ _1341_ VPWR _1342_ VGND net725 net717 sg13g2_o21ai_1
Xfanout745 net746 net745 VPWR VGND sg13g2_buf_8
Xfanout734 falu_i.falutop.alu_data_in\[11\] net734 VPWR VGND sg13g2_buf_2
Xfanout756 net757 net756 VPWR VGND sg13g2_buf_2
Xfanout767 falu_i.falutop.alu_data_in\[1\] net767 VPWR VGND sg13g2_buf_8
X_5420__212 VPWR VGND net212 sg13g2_tiehi
Xfanout789 net790 net789 VPWR VGND sg13g2_buf_8
Xfanout778 net779 net778 VPWR VGND sg13g2_buf_8
XFILLER_14_504 VPWR VGND sg13g2_fill_1
XFILLER_41_334 VPWR VGND sg13g2_fill_2
XFILLER_10_776 VPWR VGND sg13g2_fill_2
XFILLER_2_953 VPWR VGND sg13g2_decap_8
XFILLER_49_412 VPWR VGND sg13g2_decap_4
XFILLER_49_434 VPWR VGND sg13g2_decap_8
XFILLER_37_607 VPWR VGND sg13g2_fill_2
XFILLER_49_489 VPWR VGND sg13g2_decap_8
XFILLER_37_629 VPWR VGND sg13g2_decap_4
XFILLER_18_865 VPWR VGND sg13g2_decap_8
XFILLER_32_301 VPWR VGND sg13g2_decap_4
XFILLER_32_323 VPWR VGND sg13g2_decap_8
XFILLER_33_835 VPWR VGND sg13g2_fill_2
XFILLER_32_356 VPWR VGND sg13g2_fill_1
XFILLER_33_857 VPWR VGND sg13g2_decap_4
XFILLER_20_529 VPWR VGND sg13g2_fill_2
X_3760_ _0908_ ppwm_i.u_ppwm.u_mem.programming _0906_ VPWR VGND sg13g2_nand2_1
XFILLER_13_581 VPWR VGND sg13g2_decap_4
X_3691_ net577 VPWR _0853_ VGND ppwm_i.u_ppwm.pwm_value\[4\] net581 sg13g2_o21ai_1
XFILLER_9_574 VPWR VGND sg13g2_fill_2
X_5430_ net171 VGND VPWR net503 ppwm_i.u_ppwm.u_mem.memory\[89\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_5361_ net330 VGND VPWR net966 ppwm_i.u_ppwm.u_mem.memory\[20\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_2
X_5292_ net113 VGND VPWR _0054_ ppwm_i.u_ppwm.global_counter\[9\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
X_4312_ net740 _2304_ _1265_ VPWR VGND sg13g2_nor2_1
X_4243_ net396 net606 _1205_ VPWR VGND sg13g2_nor2_1
X_4174_ net819 VPWR _1152_ VGND net1037 net636 sg13g2_o21ai_1
X_3125_ _2439_ _0360_ _0361_ VPWR VGND sg13g2_nor2_1
X_3056_ _2410_ _2408_ _2409_ _2407_ _2406_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_802 VPWR VGND sg13g2_decap_8
XFILLER_23_312 VPWR VGND sg13g2_fill_1
XFILLER_24_879 VPWR VGND sg13g2_decap_8
XFILLER_11_529 VPWR VGND sg13g2_decap_8
X_3958_ VGND VPWR _2165_ net674 _0198_ _1007_ sg13g2_a21oi_1
X_3889_ net835 VPWR _0973_ VGND net522 net647 sg13g2_o21ai_1
X_2909_ VPWR _2263_ ppwm_i.u_ppwm.global_counter\[14\] VGND sg13g2_inv_1
X_5559_ net157 VGND VPWR net1154 falu_i.falutop.alu_data_in\[5\] clknet_leaf_36_clk
+ sg13g2_dfrbpq_2
Xfanout575 _0617_ net575 VPWR VGND sg13g2_buf_8
Xfanout564 net565 net564 VPWR VGND sg13g2_buf_2
Xfanout597 _2404_ net597 VPWR VGND sg13g2_buf_2
Xfanout586 _2375_ net586 VPWR VGND sg13g2_buf_8
XFILLER_19_618 VPWR VGND sg13g2_fill_1
XFILLER_19_629 VPWR VGND sg13g2_decap_4
XFILLER_14_345 VPWR VGND sg13g2_fill_1
XFILLER_15_868 VPWR VGND sg13g2_decap_8
XFILLER_41_153 VPWR VGND sg13g2_decap_4
XFILLER_41_186 VPWR VGND sg13g2_fill_1
XFILLER_6_511 VPWR VGND sg13g2_fill_2
XFILLER_2_794 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_fill_1
XFILLER_2_11 VPWR VGND sg13g2_decap_8
XFILLER_49_297 VPWR VGND sg13g2_decap_8
XFILLER_18_651 VPWR VGND sg13g2_fill_2
XFILLER_46_993 VPWR VGND sg13g2_decap_8
X_4930_ _1871_ _1870_ _1843_ _1874_ VPWR VGND sg13g2_a21o_1
XFILLER_18_695 VPWR VGND sg13g2_decap_8
X_4861_ VGND VPWR net727 _1803_ _1806_ _1802_ sg13g2_a21oi_1
XFILLER_21_805 VPWR VGND sg13g2_decap_8
XFILLER_36_1018 VPWR VGND sg13g2_decap_8
XFILLER_32_142 VPWR VGND sg13g2_fill_1
XFILLER_32_164 VPWR VGND sg13g2_fill_1
X_3812_ VGND VPWR _2216_ net655 _0125_ _0934_ sg13g2_a21oi_1
X_4792_ _1728_ _1734_ _1736_ _1737_ _1738_ VPWR VGND sg13g2_nor4_1
X_3743_ _0805_ net570 _0899_ _0900_ VPWR VGND sg13g2_nor3_1
X_3674_ VPWR VGND _0679_ net798 _0837_ _2241_ _0084_ net570 sg13g2_a221oi_1
X_5413_ net226 VGND VPWR _0172_ ppwm_i.u_ppwm.u_mem.memory\[72\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_5344_ net364 VGND VPWR net561 ppwm_i.u_ppwm.u_mem.memory\[3\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_5275_ net146 VGND VPWR _0037_ ppwm_i.u_ppwm.u_pwm.counter\[3\] clknet_leaf_14_clk
+ sg13g2_dfrbpq_2
X_4226_ VGND VPWR net780 falu_i.falutop.div_inst.a\[2\] _1192_ _1191_ sg13g2_a21oi_1
X_4157_ net1085 net983 _1103_ _0260_ VPWR VGND sg13g2_mux2_1
X_3108_ VGND VPWR net801 _0347_ _0007_ _0348_ sg13g2_a21oi_1
XFILLER_29_949 VPWR VGND sg13g2_decap_8
XFILLER_37_971 VPWR VGND sg13g2_decap_8
X_4088_ _1092_ _1048_ _1088_ VPWR VGND sg13g2_nand2_1
XFILLER_15_109 VPWR VGND sg13g2_fill_1
X_3039_ _2393_ net690 _2169_ net697 _2173_ VPWR VGND sg13g2_a22oi_1
X_5270__156 VPWR VGND net156 sg13g2_tiehi
XFILLER_20_860 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_4_1027 VPWR VGND sg13g2_fill_2
XFILLER_43_996 VPWR VGND sg13g2_decap_8
XFILLER_15_698 VPWR VGND sg13g2_fill_2
XFILLER_11_860 VPWR VGND sg13g2_decap_8
XFILLER_30_668 VPWR VGND sg13g2_fill_2
XFILLER_7_853 VPWR VGND sg13g2_decap_8
XFILLER_6_352 VPWR VGND sg13g2_decap_4
X_3390_ _0568_ net592 _0567_ VPWR VGND sg13g2_nand2b_1
XFILLER_35_4 VPWR VGND sg13g2_fill_1
X_5060_ _1986_ _2000_ _2001_ VPWR VGND sg13g2_nor2_1
XFILLER_42_1022 VPWR VGND sg13g2_decap_8
X_4011_ _1040_ net1156 _0217_ VPWR VGND sg13g2_and2_1
XFILLER_37_212 VPWR VGND sg13g2_fill_2
X_5340__371 VPWR VGND net371 sg13g2_tiehi
XFILLER_19_982 VPWR VGND sg13g2_decap_8
X_4913_ _1810_ VPWR _1857_ VGND _1752_ _1811_ sg13g2_o21ai_1
XFILLER_34_941 VPWR VGND sg13g2_decap_8
X_4844_ _1774_ VPWR _1789_ VGND _1684_ _1775_ sg13g2_o21ai_1
X_4775_ _1720_ _1719_ _1721_ VPWR VGND sg13g2_nor2b_1
XFILLER_20_145 VPWR VGND sg13g2_decap_4
X_3726_ _0882_ _0883_ _0865_ _0884_ VPWR VGND sg13g2_nand3_1
X_3657_ _0822_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] net609 VPWR VGND sg13g2_nand2_1
X_3588_ _0758_ _0757_ _0622_ _0720_ net571 VPWR VGND sg13g2_a22oi_1
X_5327_ net47 VGND VPWR _0086_ ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] clknet_leaf_13_clk
+ sg13g2_dfrbpq_2
XFILLER_0_539 VPWR VGND sg13g2_decap_8
X_5258_ net179 VGND VPWR _0020_ falu_i.falutop.i2c_inst.data_in\[16\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_4209_ _1178_ VPWR _1179_ VGND net931 net567 sg13g2_o21ai_1
X_5189_ VGND VPWR _2297_ net617 _0327_ _2109_ sg13g2_a21oi_1
XFILLER_29_735 VPWR VGND sg13g2_decap_4
XFILLER_19_1024 VPWR VGND sg13g2_decap_4
XFILLER_25_974 VPWR VGND sg13g2_decap_8
XFILLER_11_101 VPWR VGND sg13g2_fill_2
XFILLER_40_988 VPWR VGND sg13g2_decap_8
XFILLER_12_668 VPWR VGND sg13g2_decap_4
XFILLER_8_639 VPWR VGND sg13g2_decap_8
XFILLER_22_63 VPWR VGND sg13g2_decap_4
XFILLER_22_74 VPWR VGND sg13g2_decap_4
XFILLER_4_845 VPWR VGND sg13g2_decap_8
XFILLER_26_1028 VPWR VGND sg13g2_fill_1
X_5504__267 VPWR VGND net267 sg13g2_tiehi
XFILLER_47_543 VPWR VGND sg13g2_fill_1
XFILLER_34_204 VPWR VGND sg13g2_fill_2
XFILLER_35_738 VPWR VGND sg13g2_fill_2
XFILLER_16_930 VPWR VGND sg13g2_decap_8
XFILLER_34_248 VPWR VGND sg13g2_decap_8
XFILLER_31_911 VPWR VGND sg13g2_fill_1
X_2890_ net1176 _2244_ VPWR VGND sg13g2_inv_4
X_4560_ net734 net759 _1324_ _1510_ VPWR VGND sg13g2_or3_1
XFILLER_30_476 VPWR VGND sg13g2_decap_4
XFILLER_6_160 VPWR VGND sg13g2_fill_1
X_4491_ _1228_ VPWR _1442_ VGND _1304_ _1321_ sg13g2_o21ai_1
X_3511_ net573 _0680_ _0684_ _0685_ VPWR VGND sg13g2_nor3_1
X_3442_ _0618_ _2344_ _0616_ VPWR VGND sg13g2_nand2_2
X_3373_ _2238_ ppwm_i.u_ppwm.global_counter\[5\] _0551_ VPWR VGND sg13g2_nor2_1
X_5112_ _2050_ _2051_ _0308_ VPWR VGND sg13g2_nor2_1
X_5043_ _1959_ _1935_ _1961_ _1984_ VPWR VGND sg13g2_a21o_1
Xheichips25_tiny_wrapper_25 VPWR VGND uo_out[2] sg13g2_tielo
Xheichips25_tiny_wrapper_14 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_22_922 VPWR VGND sg13g2_decap_8
X_4827_ _1773_ _1748_ _1772_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_999 VPWR VGND sg13g2_decap_8
X_4758_ _1686_ _1703_ _1705_ VPWR VGND sg13g2_nor2b_1
XFILLER_49_1006 VPWR VGND sg13g2_decap_8
X_3709_ net575 VPWR _0869_ VGND _0864_ _0867_ sg13g2_o21ai_1
X_4689_ _1637_ _1620_ _1635_ VPWR VGND sg13g2_xnor2_1
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_fill_1
XFILLER_49_808 VPWR VGND sg13g2_decap_8
XFILLER_48_307 VPWR VGND sg13g2_decap_4
XFILLER_1_1008 VPWR VGND sg13g2_decap_8
XFILLER_44_568 VPWR VGND sg13g2_decap_4
XFILLER_13_922 VPWR VGND sg13g2_decap_8
XFILLER_40_741 VPWR VGND sg13g2_fill_1
XFILLER_9_937 VPWR VGND sg13g2_decap_8
XFILLER_13_999 VPWR VGND sg13g2_decap_8
XFILLER_32_1010 VPWR VGND sg13g2_decap_8
XFILLER_33_95 VPWR VGND sg13g2_fill_1
XFILLER_4_675 VPWR VGND sg13g2_decap_8
Xhold3 ppwm_i.u_ppwm.u_mem.clk_prog_sync2 VPWR VGND net375 sg13g2_dlygate4sd3_1
XFILLER_47_362 VPWR VGND sg13g2_fill_2
XFILLER_47_351 VPWR VGND sg13g2_fill_2
X_3991_ net680 VPWR _1026_ VGND net1152 net378 sg13g2_o21ai_1
X_2942_ net721 _2296_ VPWR VGND sg13g2_inv_4
XFILLER_16_771 VPWR VGND sg13g2_decap_8
XFILLER_16_782 VPWR VGND sg13g2_fill_1
X_2873_ VPWR _2227_ net888 VGND sg13g2_inv_1
X_4612_ _1559_ _1560_ _1561_ VPWR VGND sg13g2_nor2_1
X_4543_ _1492_ _1482_ _1493_ VPWR VGND sg13g2_xor2_1
Xhold425 _0063_ VPWR VGND net1077 sg13g2_dlygate4sd3_1
Xhold414 ppwm_i.u_ppwm.u_pwm.counter\[6\] VPWR VGND net1066 sg13g2_dlygate4sd3_1
Xhold436 falu_i.falutop.i2c_inst.result\[6\] VPWR VGND net1088 sg13g2_dlygate4sd3_1
Xhold403 _0262_ VPWR VGND net1055 sg13g2_dlygate4sd3_1
Xhold447 _0273_ VPWR VGND net1099 sg13g2_dlygate4sd3_1
X_4474_ VGND VPWR _1425_ _1424_ _1399_ sg13g2_or2_1
Xhold458 falu_i.falutop.div_inst.rem\[2\] VPWR VGND net1110 sg13g2_dlygate4sd3_1
Xhold469 _0442_ VPWR VGND net1121 sg13g2_dlygate4sd3_1
X_5407__238 VPWR VGND net238 sg13g2_tiehi
X_3425_ _0603_ _2419_ _0602_ VPWR VGND sg13g2_nand2_1
X_3356_ _0534_ ppwm_i.u_ppwm.global_counter\[1\] net784 VPWR VGND sg13g2_nand2b_1
X_3287_ _0469_ VPWR _0470_ VGND _2275_ ppwm_i.u_ppwm.u_pwm.cmp_value\[6\] sg13g2_o21ai_1
X_5381__290 VPWR VGND net290 sg13g2_tiehi
X_5522__186 VPWR VGND net186 sg13g2_tiehi
X_5026_ _1968_ net615 _1966_ _1967_ VPWR VGND sg13g2_and3_2
XFILLER_38_373 VPWR VGND sg13g2_decap_8
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_13_218 VPWR VGND sg13g2_fill_1
XFILLER_10_936 VPWR VGND sg13g2_decap_8
X_5539__68 VPWR VGND net68 sg13g2_tiehi
XFILLER_22_796 VPWR VGND sg13g2_decap_8
X_5464__365 VPWR VGND net365 sg13g2_tiehi
XFILLER_0_122 VPWR VGND sg13g2_decap_8
XFILLER_1_656 VPWR VGND sg13g2_fill_2
XFILLER_0_166 VPWR VGND sg13g2_fill_2
XFILLER_29_351 VPWR VGND sg13g2_decap_8
XFILLER_29_362 VPWR VGND sg13g2_fill_2
XFILLER_28_95 VPWR VGND sg13g2_fill_2
XFILLER_9_734 VPWR VGND sg13g2_decap_8
XFILLER_40_593 VPWR VGND sg13g2_decap_8
XFILLER_9_789 VPWR VGND sg13g2_decap_4
XFILLER_5_951 VPWR VGND sg13g2_decap_8
XFILLER_4_450 VPWR VGND sg13g2_decap_8
X_3210_ _0417_ net1177 _0415_ VPWR VGND sg13g2_nand2_1
X_4190_ net803 VPWR _1164_ VGND net1110 net634 sg13g2_o21ai_1
X_3141_ _2446_ net1007 _0372_ VPWR VGND sg13g2_nor2_1
X_3072_ _2424_ net981 net821 _0000_ VPWR VGND sg13g2_nand3_1
XFILLER_35_354 VPWR VGND sg13g2_fill_1
XFILLER_23_549 VPWR VGND sg13g2_fill_1
X_3974_ VGND VPWR _2159_ net672 _0206_ _1015_ sg13g2_a21oi_1
X_2925_ VPWR _2279_ net535 VGND sg13g2_inv_1
X_2856_ VPWR _2210_ net472 VGND sg13g2_inv_1
Xhold211 ppwm_i.u_ppwm.u_pwm.counter\[3\] VPWR VGND net863 sg13g2_dlygate4sd3_1
X_5575_ net359 VGND VPWR net984 falu_i.falutop.div_inst.b\[5\] clknet_leaf_4_clk sg13g2_dfrbpq_1
Xhold200 ppwm_i.u_ppwm.u_mem.memory\[3\] VPWR VGND net852 sg13g2_dlygate4sd3_1
Xhold233 ppwm_i.u_ppwm.u_mem.memory\[60\] VPWR VGND net885 sg13g2_dlygate4sd3_1
X_4526_ _1476_ _1463_ _1474_ VPWR VGND sg13g2_xnor2_1
Xhold222 _0236_ VPWR VGND net874 sg13g2_dlygate4sd3_1
Xhold244 ppwm_i.u_ppwm.u_mem.memory\[12\] VPWR VGND net896 sg13g2_dlygate4sd3_1
Xhold255 _0336_ VPWR VGND net907 sg13g2_dlygate4sd3_1
Xhold266 _1142_ VPWR VGND net918 sg13g2_dlygate4sd3_1
X_4457_ _1403_ _1408_ _0296_ VPWR VGND sg13g2_nor2_1
Xhold277 _0113_ VPWR VGND net929 sg13g2_dlygate4sd3_1
X_3408_ _0586_ _2258_ net591 VPWR VGND sg13g2_nand2_1
Xfanout713 net714 net713 VPWR VGND sg13g2_buf_1
Xhold288 _1147_ VPWR VGND net940 sg13g2_dlygate4sd3_1
Xfanout724 falu_i.falutop.alu_data_in\[13\] net724 VPWR VGND sg13g2_buf_8
Xhold299 ppwm_i.u_ppwm.u_mem.memory\[111\] VPWR VGND net951 sg13g2_dlygate4sd3_1
Xfanout702 net703 net702 VPWR VGND sg13g2_buf_8
X_4388_ net710 _1293_ _1341_ VPWR VGND sg13g2_nor2_1
Xfanout746 falu_i.falutop.alu_data_in\[8\] net746 VPWR VGND sg13g2_buf_8
Xfanout757 net758 net757 VPWR VGND sg13g2_buf_1
Xfanout735 net736 net735 VPWR VGND sg13g2_buf_8
X_3339_ _0517_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] _2243_ VPWR VGND sg13g2_nand2_1
Xfanout779 net887 net779 VPWR VGND sg13g2_buf_8
Xfanout768 net769 net768 VPWR VGND sg13g2_buf_8
XFILLER_22_1020 VPWR VGND sg13g2_decap_8
X_5009_ _1951_ net718 net751 VPWR VGND sg13g2_nand2_1
XFILLER_14_516 VPWR VGND sg13g2_decap_4
XFILLER_14_538 VPWR VGND sg13g2_decap_8
XFILLER_10_700 VPWR VGND sg13g2_decap_4
XFILLER_22_571 VPWR VGND sg13g2_decap_4
XFILLER_10_744 VPWR VGND sg13g2_decap_4
XFILLER_14_64 VPWR VGND sg13g2_fill_2
XFILLER_2_932 VPWR VGND sg13g2_decap_8
X_5280__136 VPWR VGND net136 sg13g2_tiehi
XFILLER_7_1014 VPWR VGND sg13g2_decap_8
XFILLER_36_107 VPWR VGND sg13g2_decap_4
XFILLER_17_321 VPWR VGND sg13g2_fill_2
XFILLER_18_844 VPWR VGND sg13g2_decap_8
XFILLER_32_379 VPWR VGND sg13g2_fill_2
XFILLER_9_564 VPWR VGND sg13g2_decap_4
X_3690_ _0851_ VPWR _0852_ VGND _0848_ _0849_ sg13g2_o21ai_1
X_5360_ net332 VGND VPWR net876 ppwm_i.u_ppwm.u_mem.memory\[19\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_5291_ net115 VGND VPWR net555 ppwm_i.u_ppwm.global_counter\[8\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
X_4311_ _1264_ net764 net739 VPWR VGND sg13g2_nand2b_1
XFILLER_45_1020 VPWR VGND sg13g2_decap_8
X_5541__52 VPWR VGND net52 sg13g2_tiehi
X_4242_ VGND VPWR net780 falu_i.falutop.div_inst.a\[6\] _1204_ _1203_ sg13g2_a21oi_1
X_4173_ VGND VPWR _2148_ net636 _0269_ _1151_ sg13g2_a21oi_1
X_3124_ _0360_ _2154_ net1017 VPWR VGND sg13g2_nand2_2
X_3055_ VPWR VGND _2183_ net790 net695 _2177_ _2409_ net703 sg13g2_a221oi_1
X_5554__219 VPWR VGND net219 sg13g2_tiehi
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_24_858 VPWR VGND sg13g2_decap_8
XFILLER_11_519 VPWR VGND sg13g2_fill_2
X_3957_ net837 VPWR _1007_ VGND net562 net674 sg13g2_o21ai_1
X_2908_ _2262_ net1180 VPWR VGND sg13g2_inv_2
X_3888_ VGND VPWR _2190_ net671 _0163_ _0972_ sg13g2_a21oi_1
X_2839_ VPWR _2193_ net885 VGND sg13g2_inv_1
X_5558_ net194 VGND VPWR net1115 falu_i.falutop.alu_data_in\[4\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_4509_ VGND VPWR net978 _1458_ _1460_ _1406_ sg13g2_a21oi_1
XFILLER_4_8 VPWR VGND sg13g2_decap_8
X_5489_ net303 VGND VPWR _0248_ falu_i.falutop.alu_inst.op\[0\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_2
Xfanout565 _1278_ net565 VPWR VGND sg13g2_buf_2
XFILLER_47_939 VPWR VGND sg13g2_decap_8
Xfanout598 net599 net598 VPWR VGND sg13g2_buf_8
Xfanout587 _1295_ net587 VPWR VGND sg13g2_buf_8
XFILLER_19_608 VPWR VGND sg13g2_fill_1
Xfanout576 _0617_ net576 VPWR VGND sg13g2_buf_2
Xclkbuf_leaf_38_clk clknet_3_1__leaf_clk clknet_leaf_38_clk VPWR VGND sg13g2_buf_8
XFILLER_27_696 VPWR VGND sg13g2_fill_2
XFILLER_15_847 VPWR VGND sg13g2_decap_8
XFILLER_42_699 VPWR VGND sg13g2_fill_2
XFILLER_41_165 VPWR VGND sg13g2_fill_1
XFILLER_23_891 VPWR VGND sg13g2_decap_8
XFILLER_29_1026 VPWR VGND sg13g2_fill_2
XFILLER_38_939 VPWR VGND sg13g2_decap_8
XFILLER_49_276 VPWR VGND sg13g2_decap_8
X_5477__331 VPWR VGND net331 sg13g2_tiehi
XFILLER_46_972 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk clknet_leaf_29_clk VPWR VGND sg13g2_buf_8
XFILLER_45_482 VPWR VGND sg13g2_fill_1
X_4860_ _1805_ net727 _1803_ VPWR VGND sg13g2_nand2_1
XFILLER_32_121 VPWR VGND sg13g2_fill_2
XFILLER_20_305 VPWR VGND sg13g2_fill_2
X_3811_ net824 VPWR _0934_ VGND ppwm_i.u_ppwm.u_mem.memory\[25\] net653 sg13g2_o21ai_1
X_4791_ _1280_ _1327_ _1241_ _1737_ VPWR VGND sg13g2_mux2_1
XFILLER_14_880 VPWR VGND sg13g2_decap_8
X_3742_ VGND VPWR net583 _0806_ _0899_ _0898_ sg13g2_a21oi_1
XFILLER_20_349 VPWR VGND sg13g2_decap_4
X_3673_ _0680_ net570 _0834_ _0836_ _0837_ VPWR VGND sg13g2_nor4_1
X_5412_ net228 VGND VPWR _0171_ ppwm_i.u_ppwm.u_mem.memory\[71\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_1
X_5343_ net366 VGND VPWR net853 ppwm_i.u_ppwm.u_mem.memory\[2\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
X_5274_ net148 VGND VPWR _0036_ ppwm_i.u_ppwm.u_pwm.counter\[2\] clknet_leaf_12_clk
+ sg13g2_dfrbpq_2
X_4225_ net780 _2150_ _1191_ VPWR VGND sg13g2_nor2_1
X_4156_ net1078 net999 _1103_ _0259_ VPWR VGND sg13g2_mux2_1
XFILLER_29_928 VPWR VGND sg13g2_decap_8
X_3107_ net823 VPWR _0348_ VGND net992 _0347_ sg13g2_o21ai_1
XFILLER_44_909 VPWR VGND sg13g2_decap_8
XFILLER_37_950 VPWR VGND sg13g2_decap_8
X_4087_ _1091_ _1089_ _1090_ VPWR VGND sg13g2_nand2_1
XFILLER_24_600 VPWR VGND sg13g2_decap_8
X_3038_ VGND VPWR _2164_ net694 _2392_ net709 sg13g2_a21oi_1
XFILLER_23_121 VPWR VGND sg13g2_fill_1
X_4989_ net818 VPWR _1932_ VGND net1062 net629 sg13g2_o21ai_1
XFILLER_12_839 VPWR VGND sg13g2_decap_8
XFILLER_23_187 VPWR VGND sg13g2_fill_2
XFILLER_4_1006 VPWR VGND sg13g2_decap_8
XFILLER_46_202 VPWR VGND sg13g2_fill_1
XFILLER_46_246 VPWR VGND sg13g2_decap_4
XFILLER_28_994 VPWR VGND sg13g2_decap_8
XFILLER_43_975 VPWR VGND sg13g2_decap_8
XFILLER_14_143 VPWR VGND sg13g2_decap_8
XFILLER_14_154 VPWR VGND sg13g2_fill_2
XFILLER_30_603 VPWR VGND sg13g2_fill_1
XFILLER_6_375 VPWR VGND sg13g2_fill_1
XFILLER_42_1001 VPWR VGND sg13g2_decap_8
X_4010_ _1041_ _1036_ net1155 VPWR VGND sg13g2_nand2b_1
XFILLER_28_4 VPWR VGND sg13g2_decap_4
XFILLER_38_747 VPWR VGND sg13g2_fill_1
XFILLER_19_961 VPWR VGND sg13g2_decap_8
XFILLER_26_909 VPWR VGND sg13g2_decap_8
X_4912_ _1856_ _1853_ _1855_ VPWR VGND sg13g2_xnor2_1
XFILLER_18_493 VPWR VGND sg13g2_decap_4
XFILLER_34_997 VPWR VGND sg13g2_decap_8
X_4843_ _1777_ VPWR _1788_ VGND _1739_ _1778_ sg13g2_o21ai_1
XFILLER_20_113 VPWR VGND sg13g2_fill_1
X_4774_ _1720_ net705 _1654_ VPWR VGND sg13g2_xnor2_1
XFILLER_20_135 VPWR VGND sg13g2_fill_1
X_3725_ net601 VPWR _0883_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] ppwm_i.u_ppwm.u_ex.reg_value_q\[6\]
+ sg13g2_o21ai_1
Xclkbuf_leaf_9_clk clknet_3_2__leaf_clk clknet_leaf_9_clk VPWR VGND sg13g2_buf_8
X_3656_ net799 _0821_ _0082_ VPWR VGND sg13g2_nor2_1
X_3587_ net609 _0738_ _0757_ VPWR VGND sg13g2_nor2_1
XFILLER_0_518 VPWR VGND sg13g2_decap_8
X_5326_ net49 VGND VPWR _0085_ ppwm_i.u_ppwm.u_ex.reg_value_q\[3\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_5257_ net181 VGND VPWR _0019_ falu_i.falutop.i2c_inst.data_in\[15\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_4208_ _1178_ net567 _1177_ VPWR VGND sg13g2_nand2_1
X_5188_ net1105 net617 _2109_ VPWR VGND sg13g2_nor2_1
XFILLER_29_747 VPWR VGND sg13g2_fill_1
X_4139_ VPWR _0249_ net1027 VGND sg13g2_inv_1
XFILLER_44_717 VPWR VGND sg13g2_fill_1
XFILLER_37_780 VPWR VGND sg13g2_fill_2
X_5417__218 VPWR VGND net218 sg13g2_tiehi
XFILLER_25_953 VPWR VGND sg13g2_decap_8
XFILLER_19_1003 VPWR VGND sg13g2_decap_8
XFILLER_24_452 VPWR VGND sg13g2_decap_8
X_5391__270 VPWR VGND net270 sg13g2_tiehi
XFILLER_40_967 VPWR VGND sg13g2_decap_8
XFILLER_20_691 VPWR VGND sg13g2_decap_8
XFILLER_22_97 VPWR VGND sg13g2_fill_2
XFILLER_26_1007 VPWR VGND sg13g2_decap_8
XFILLER_19_257 VPWR VGND sg13g2_fill_2
XFILLER_19_268 VPWR VGND sg13g2_fill_2
XFILLER_16_986 VPWR VGND sg13g2_decap_8
XFILLER_30_411 VPWR VGND sg13g2_decap_4
Xclkbuf_3_4__f_clk clknet_0_clk clknet_3_4__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_31_989 VPWR VGND sg13g2_decap_8
XFILLER_8_99 VPWR VGND sg13g2_fill_2
XFILLER_8_88 VPWR VGND sg13g2_decap_8
X_3510_ VGND VPWR net588 _0682_ _0684_ _0683_ sg13g2_a21oi_1
X_5327__47 VPWR VGND net47 sg13g2_tiehi
X_4490_ net631 _1440_ _1268_ _1441_ VPWR VGND sg13g2_nand3_1
X_3441_ _2344_ _0616_ _0617_ VPWR VGND sg13g2_and2_1
X_3372_ _0550_ _2237_ ppwm_i.u_ppwm.global_counter\[6\] VPWR VGND sg13g2_nand2_1
X_5111_ net815 VPWR _2051_ VGND net1035 net627 sg13g2_o21ai_1
X_5042_ VPWR VGND _1981_ _1982_ _1978_ _1933_ _1983_ _1962_ sg13g2_a221oi_1
XFILLER_38_544 VPWR VGND sg13g2_fill_1
Xheichips25_tiny_wrapper_26 VPWR VGND uo_out[3] sg13g2_tielo
Xheichips25_tiny_wrapper_15 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_19_780 VPWR VGND sg13g2_fill_2
XFILLER_22_901 VPWR VGND sg13g2_decap_8
XFILLER_21_411 VPWR VGND sg13g2_fill_2
X_4826_ _1772_ _1749_ _1769_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_978 VPWR VGND sg13g2_decap_8
XFILLER_33_282 VPWR VGND sg13g2_decap_8
X_4757_ _1704_ _1686_ _1703_ VPWR VGND sg13g2_nand2b_1
X_3708_ _0864_ _0867_ _0868_ VPWR VGND sg13g2_and2_1
X_4688_ _1636_ _1620_ _1635_ VPWR VGND sg13g2_nand2_1
X_3639_ _0586_ VPWR _0806_ VGND ppwm_i.u_ppwm.global_counter\[9\] net592 sg13g2_o21ai_1
XFILLER_1_805 VPWR VGND sg13g2_decap_8
X_5309_ net83 VGND VPWR _0068_ ppwm_i.u_ppwm.pc\[2\] clknet_leaf_22_clk sg13g2_dfrbpq_1
X_5423__200 VPWR VGND net200 sg13g2_tiehi
XFILLER_0_326 VPWR VGND sg13g2_fill_2
XFILLER_0_359 VPWR VGND sg13g2_fill_2
XFILLER_0_348 VPWR VGND sg13g2_decap_8
XFILLER_29_500 VPWR VGND sg13g2_fill_1
XFILLER_44_536 VPWR VGND sg13g2_fill_2
XFILLER_17_739 VPWR VGND sg13g2_fill_1
XFILLER_13_901 VPWR VGND sg13g2_decap_8
XFILLER_9_916 VPWR VGND sg13g2_decap_8
XFILLER_12_422 VPWR VGND sg13g2_decap_4
XFILLER_12_455 VPWR VGND sg13g2_fill_2
XFILLER_13_978 VPWR VGND sg13g2_decap_8
XFILLER_40_786 VPWR VGND sg13g2_decap_8
XFILLER_12_477 VPWR VGND sg13g2_decap_4
XFILLER_4_665 VPWR VGND sg13g2_fill_2
XFILLER_4_654 VPWR VGND sg13g2_fill_2
Xhold4 ppwm_i.u_ppwm.polarity VPWR VGND net376 sg13g2_dlygate4sd3_1
XFILLER_48_886 VPWR VGND sg13g2_decap_8
XFILLER_35_514 VPWR VGND sg13g2_fill_2
X_3990_ net1152 net378 _1025_ VPWR VGND sg13g2_and2_1
X_2941_ _2295_ net740 VPWR VGND sg13g2_inv_2
X_4611_ VGND VPWR _1557_ _1558_ _1560_ _1553_ sg13g2_a21oi_1
X_2872_ VPWR _2226_ net896 VGND sg13g2_inv_1
XFILLER_8_993 VPWR VGND sg13g2_decap_8
X_4542_ _1489_ _1491_ _1492_ VPWR VGND sg13g2_nor2_1
Xhold415 _0414_ VPWR VGND net1067 sg13g2_dlygate4sd3_1
X_4473_ _1424_ _1397_ _1422_ VPWR VGND sg13g2_xnor2_1
Xhold426 falu_i.falutop.div_inst.b1\[4\] VPWR VGND net1078 sg13g2_dlygate4sd3_1
Xhold404 falu_i.falutop.div_inst.b1\[6\] VPWR VGND net1056 sg13g2_dlygate4sd3_1
X_3424_ _0588_ _0601_ net610 _0602_ VPWR VGND sg13g2_nand3_1
Xhold448 falu_i.falutop.div_inst.rem\[6\] VPWR VGND net1100 sg13g2_dlygate4sd3_1
Xhold437 falu_i.falutop.i2c_inst.result\[3\] VPWR VGND net1089 sg13g2_dlygate4sd3_1
Xhold459 ppwm_i.u_ppwm.u_pwm.counter\[0\] VPWR VGND net1111 sg13g2_dlygate4sd3_1
X_3355_ ppwm_i.u_ppwm.pwm_value\[7\] _2268_ _0533_ VPWR VGND sg13g2_nor2_1
X_3286_ _0469_ _0467_ _0468_ _2281_ ppwm_i.u_ppwm.u_pwm.counter\[7\] VPWR VGND sg13g2_a22oi_1
XFILLER_39_853 VPWR VGND sg13g2_decap_8
X_5025_ _1919_ _1921_ _1965_ _1967_ VPWR VGND sg13g2_or3_1
XFILLER_39_864 VPWR VGND sg13g2_fill_1
XFILLER_38_385 VPWR VGND sg13g2_decap_4
XFILLER_26_525 VPWR VGND sg13g2_fill_1
X_5492__297 VPWR VGND net297 sg13g2_tiehi
XFILLER_34_580 VPWR VGND sg13g2_fill_1
XFILLER_10_915 VPWR VGND sg13g2_decap_8
XFILLER_16_1028 VPWR VGND sg13g2_fill_1
XFILLER_22_775 VPWR VGND sg13g2_decap_8
X_4809_ _1755_ net766 net719 net768 net713 VPWR VGND sg13g2_a22oi_1
XFILLER_1_635 VPWR VGND sg13g2_fill_1
XFILLER_45_801 VPWR VGND sg13g2_fill_2
XFILLER_17_547 VPWR VGND sg13g2_fill_2
XFILLER_45_867 VPWR VGND sg13g2_fill_1
XFILLER_44_333 VPWR VGND sg13g2_fill_2
XFILLER_17_569 VPWR VGND sg13g2_decap_8
XFILLER_13_720 VPWR VGND sg13g2_decap_8
XFILLER_9_702 VPWR VGND sg13g2_decap_8
XFILLER_9_713 VPWR VGND sg13g2_fill_2
XFILLER_9_757 VPWR VGND sg13g2_decap_8
XFILLER_5_930 VPWR VGND sg13g2_decap_8
X_3140_ VGND VPWR net800 _0370_ _0016_ _0371_ sg13g2_a21oi_1
XFILLER_10_4 VPWR VGND sg13g2_fill_2
X_3071_ _2425_ net980 ppwm_i.u_ppwm.period_start VPWR VGND sg13g2_nand2b_1
XFILLER_35_311 VPWR VGND sg13g2_fill_1
XFILLER_35_344 VPWR VGND sg13g2_fill_2
X_3973_ net837 VPWR _1015_ VGND ppwm_i.u_ppwm.u_mem.memory\[106\] net672 sg13g2_o21ai_1
X_2924_ VPWR _2278_ net863 VGND sg13g2_inv_1
X_2855_ VPWR _2209_ net424 VGND sg13g2_inv_1
X_5241__93 VPWR VGND net93 sg13g2_tiehi
X_5574_ net367 VGND VPWR net1000 falu_i.falutop.div_inst.b\[4\] clknet_leaf_3_clk
+ sg13g2_dfrbpq_1
X_4525_ _1475_ _1463_ _1474_ VPWR VGND sg13g2_nand2_1
Xhold201 _0102_ VPWR VGND net853 sg13g2_dlygate4sd3_1
Xhold234 ppwm_i.u_ppwm.u_mem.memory\[80\] VPWR VGND net886 sg13g2_dlygate4sd3_1
Xhold212 _0406_ VPWR VGND net864 sg13g2_dlygate4sd3_1
Xhold223 ppwm_i.u_ppwm.u_mem.memory\[19\] VPWR VGND net875 sg13g2_dlygate4sd3_1
Xhold245 ppwm_i.u_ppwm.u_mem.memory\[34\] VPWR VGND net897 sg13g2_dlygate4sd3_1
Xhold278 ppwm_i.u_ppwm.u_mem.memory\[83\] VPWR VGND net930 sg13g2_dlygate4sd3_1
X_4456_ _1402_ VPWR _1408_ VGND _1406_ _1407_ sg13g2_o21ai_1
Xhold267 _0253_ VPWR VGND net919 sg13g2_dlygate4sd3_1
Xhold256 falu_i.falutop.i2c_inst.data_in\[15\] VPWR VGND net908 sg13g2_dlygate4sd3_1
X_3407_ ppwm_i.u_ppwm.global_counter\[18\] _0581_ _0585_ VPWR VGND net782 sg13g2_nand3b_1
Xhold289 _0265_ VPWR VGND net941 sg13g2_dlygate4sd3_1
Xfanout714 net715 net714 VPWR VGND sg13g2_buf_8
X_4387_ _1340_ _1289_ _1339_ VPWR VGND sg13g2_nand2b_1
Xfanout703 net704 net703 VPWR VGND sg13g2_buf_8
X_3338_ _2330_ _2344_ net419 _0516_ VPWR VGND _2360_ sg13g2_nand4_1
Xfanout747 net748 net747 VPWR VGND sg13g2_buf_8
Xfanout725 net726 net725 VPWR VGND sg13g2_buf_8
Xfanout758 net759 net758 VPWR VGND sg13g2_buf_1
Xfanout736 net739 net736 VPWR VGND sg13g2_buf_8
Xfanout769 net770 net769 VPWR VGND sg13g2_buf_8
X_3269_ ppwm_i.u_ppwm.global_counter\[16\] _0452_ net989 _0455_ VPWR VGND sg13g2_nand3_1
XFILLER_46_609 VPWR VGND sg13g2_decap_8
XFILLER_45_119 VPWR VGND sg13g2_fill_2
X_5008_ _1803_ _1949_ _1950_ VPWR VGND sg13g2_nor2_1
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_2_911 VPWR VGND sg13g2_decap_8
XFILLER_2_988 VPWR VGND sg13g2_decap_8
XFILLER_39_62 VPWR VGND sg13g2_fill_2
XFILLER_49_469 VPWR VGND sg13g2_fill_2
XFILLER_39_95 VPWR VGND sg13g2_fill_2
XFILLER_18_823 VPWR VGND sg13g2_decap_8
XFILLER_44_185 VPWR VGND sg13g2_fill_2
XFILLER_32_347 VPWR VGND sg13g2_decap_8
X_5290_ net117 VGND VPWR _0052_ ppwm_i.u_ppwm.global_counter\[7\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_2
X_4310_ _1263_ net759 net734 VPWR VGND sg13g2_nand2b_1
X_4241_ net780 _2146_ _1203_ VPWR VGND sg13g2_nor2_1
X_4172_ net818 VPWR _1151_ VGND net937 net636 sg13g2_o21ai_1
X_3123_ net1016 falu_i.falutop.i2c_inst.counter\[3\] _0359_ VPWR VGND sg13g2_nor2b_2
XFILLER_49_992 VPWR VGND sg13g2_decap_8
X_3054_ _2408_ net691 _2188_ net697 _2193_ VPWR VGND sg13g2_a22oi_1
XFILLER_24_837 VPWR VGND sg13g2_decap_8
X_3956_ VGND VPWR _2166_ net674 _0197_ _1006_ sg13g2_a21oi_1
X_2907_ VPWR _2261_ ppwm_i.u_ppwm.global_counter\[16\] VGND sg13g2_inv_1
X_3887_ net835 VPWR _0972_ VGND ppwm_i.u_ppwm.u_mem.memory\[63\] net671 sg13g2_o21ai_1
X_5350__352 VPWR VGND net352 sg13g2_tiehi
X_2838_ VPWR _2192_ net437 VGND sg13g2_inv_1
X_5557_ net202 VGND VPWR net1136 falu_i.falutop.alu_data_in\[3\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_4508_ VGND VPWR _1459_ _1458_ net978 sg13g2_or2_1
X_5488_ net305 VGND VPWR _0247_ falu_i.falutop.div_inst.done clknet_leaf_44_clk sg13g2_dfrbpq_2
X_4439_ _1372_ _1377_ _1386_ _1390_ _1391_ VPWR VGND sg13g2_nor4_1
Xfanout566 _1278_ net566 VPWR VGND sg13g2_buf_8
XFILLER_47_918 VPWR VGND sg13g2_decap_8
Xfanout577 net580 net577 VPWR VGND sg13g2_buf_8
Xfanout599 _2404_ net599 VPWR VGND sg13g2_buf_8
Xfanout588 net590 net588 VPWR VGND sg13g2_buf_8
XFILLER_46_439 VPWR VGND sg13g2_decap_8
XFILLER_27_631 VPWR VGND sg13g2_fill_1
XFILLER_15_826 VPWR VGND sg13g2_decap_8
XFILLER_26_174 VPWR VGND sg13g2_decap_8
XFILLER_23_870 VPWR VGND sg13g2_decap_8
XFILLER_6_502 VPWR VGND sg13g2_fill_1
XFILLER_22_391 VPWR VGND sg13g2_decap_4
XFILLER_6_535 VPWR VGND sg13g2_decap_8
XFILLER_6_546 VPWR VGND sg13g2_fill_2
XFILLER_29_1005 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_fill_1
XFILLER_2_763 VPWR VGND sg13g2_fill_2
XFILLER_49_244 VPWR VGND sg13g2_decap_8
XFILLER_38_929 VPWR VGND sg13g2_decap_4
XFILLER_46_951 VPWR VGND sg13g2_decap_8
XFILLER_17_141 VPWR VGND sg13g2_fill_2
XFILLER_17_152 VPWR VGND sg13g2_fill_2
XFILLER_32_100 VPWR VGND sg13g2_fill_1
X_4790_ VGND VPWR _1242_ _1323_ _1736_ _1735_ sg13g2_a21oi_1
X_3810_ VGND VPWR _2217_ net659 _0124_ _0933_ sg13g2_a21oi_1
X_3741_ net580 VPWR _0898_ VGND ppwm_i.u_ppwm.pwm_value\[9\] net583 sg13g2_o21ai_1
X_5256__183 VPWR VGND net183 sg13g2_tiehi
XFILLER_20_317 VPWR VGND sg13g2_decap_8
X_3672_ VGND VPWR net582 _0682_ _0836_ _0835_ sg13g2_a21oi_1
X_5411_ net230 VGND VPWR net416 ppwm_i.u_ppwm.u_mem.memory\[70\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_5342_ net368 VGND VPWR net524 ppwm_i.u_ppwm.u_mem.memory\[1\] clknet_leaf_33_clk
+ sg13g2_dfrbpq_1
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_5_590 VPWR VGND sg13g2_decap_8
X_5273_ net150 VGND VPWR _0035_ ppwm_i.u_ppwm.u_pwm.counter\[1\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
X_4224_ VGND VPWR net605 _1189_ _0281_ _1190_ sg13g2_a21oi_1
X_4155_ VPWR _0258_ net995 VGND sg13g2_inv_1
X_3106_ _2434_ net1014 _0347_ VPWR VGND sg13g2_nor2_1
X_4086_ _1090_ _0343_ falu_i.falutop.i2c_inst.result\[6\] _2445_ falu_i.falutop.i2c_inst.result\[5\]
+ VPWR VGND sg13g2_a22oi_1
X_5378__296 VPWR VGND net296 sg13g2_tiehi
X_3037_ _2391_ net702 ppwm_i.u_ppwm.u_mem.memory\[108\] VPWR VGND sg13g2_nand2b_1
XFILLER_36_450 VPWR VGND sg13g2_decap_8
XFILLER_36_472 VPWR VGND sg13g2_fill_2
XFILLER_24_645 VPWR VGND sg13g2_fill_1
XFILLER_24_678 VPWR VGND sg13g2_fill_1
X_4988_ VPWR VGND net638 net630 _1930_ net614 _1931_ _1927_ sg13g2_a221oi_1
X_3939_ net836 VPWR _0998_ VGND ppwm_i.u_ppwm.u_mem.memory\[90\] net646 sg13g2_o21ai_1
XFILLER_20_895 VPWR VGND sg13g2_decap_8
XFILLER_3_549 VPWR VGND sg13g2_fill_2
XFILLER_47_704 VPWR VGND sg13g2_fill_2
XFILLER_27_461 VPWR VGND sg13g2_fill_2
XFILLER_28_973 VPWR VGND sg13g2_decap_8
XFILLER_36_63 VPWR VGND sg13g2_fill_1
XFILLER_43_954 VPWR VGND sg13g2_decap_8
XFILLER_27_494 VPWR VGND sg13g2_fill_2
XFILLER_42_464 VPWR VGND sg13g2_fill_1
XFILLER_15_667 VPWR VGND sg13g2_decap_8
XFILLER_42_497 VPWR VGND sg13g2_decap_8
XFILLER_7_800 VPWR VGND sg13g2_decap_8
XFILLER_11_895 VPWR VGND sg13g2_decap_8
XFILLER_7_888 VPWR VGND sg13g2_decap_8
XFILLER_2_582 VPWR VGND sg13g2_fill_1
XFILLER_38_704 VPWR VGND sg13g2_fill_2
XFILLER_19_940 VPWR VGND sg13g2_decap_8
XFILLER_46_792 VPWR VGND sg13g2_fill_1
X_4911_ _1855_ _1622_ _1753_ VPWR VGND sg13g2_xnor2_1
XFILLER_33_464 VPWR VGND sg13g2_fill_1
XFILLER_34_976 VPWR VGND sg13g2_decap_8
X_4842_ _1309_ VPWR _1787_ VGND _1721_ _1786_ sg13g2_o21ai_1
XFILLER_33_497 VPWR VGND sg13g2_decap_4
X_4773_ _1657_ VPWR _1719_ VGND _1595_ _1655_ sg13g2_o21ai_1
X_3724_ _0856_ _0864_ _0850_ _0882_ VPWR VGND _0874_ sg13g2_nand4_1
X_3655_ _0820_ VPWR _0821_ VGND net1173 _0813_ sg13g2_o21ai_1
X_3586_ _0755_ VPWR _0756_ VGND _0627_ _0714_ sg13g2_o21ai_1
X_5325_ net51 VGND VPWR _0084_ ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_5525__174 VPWR VGND net174 sg13g2_tiehi
X_5256_ net183 VGND VPWR _0018_ falu_i.falutop.i2c_inst.data_in\[14\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_4207_ _1177_ _1127_ _1128_ VPWR VGND sg13g2_xnor2_1
X_5187_ VGND VPWR _2296_ net617 _0326_ _2108_ sg13g2_a21oi_1
X_4138_ _1137_ falu_i.falutop.alu_inst.op\[1\] net619 net833 net1026 VPWR VGND sg13g2_a22oi_1
XFILLER_28_247 VPWR VGND sg13g2_decap_4
XFILLER_43_206 VPWR VGND sg13g2_fill_2
X_4069_ net945 falu_i.falutop.data_in\[10\] net685 _0238_ VPWR VGND sg13g2_mux2_1
XFILLER_25_932 VPWR VGND sg13g2_decap_8
XFILLER_40_946 VPWR VGND sg13g2_decap_8
XFILLER_8_619 VPWR VGND sg13g2_fill_2
X_5467__353 VPWR VGND net353 sg13g2_tiehi
XFILLER_34_228 VPWR VGND sg13g2_fill_1
XFILLER_43_762 VPWR VGND sg13g2_fill_1
XFILLER_16_965 VPWR VGND sg13g2_decap_8
XFILLER_27_291 VPWR VGND sg13g2_fill_2
XFILLER_15_464 VPWR VGND sg13g2_decap_4
XFILLER_30_456 VPWR VGND sg13g2_decap_8
XFILLER_31_968 VPWR VGND sg13g2_decap_8
XFILLER_11_692 VPWR VGND sg13g2_fill_2
X_3440_ _2329_ _2360_ _0616_ VPWR VGND sg13g2_nor2_2
X_3371_ VGND VPWR _2243_ ppwm_i.u_ppwm.global_counter\[9\] _0549_ net591 sg13g2_a21oi_1
X_5110_ VPWR VGND net638 net630 _2049_ net614 _2050_ _2046_ sg13g2_a221oi_1
X_5041_ _1963_ _1919_ _1982_ VPWR VGND sg13g2_nor2b_1
XFILLER_38_512 VPWR VGND sg13g2_fill_1
Xheichips25_tiny_wrapper_16 VPWR VGND uio_out[0] sg13g2_tielo
Xheichips25_tiny_wrapper_27 VPWR VGND uo_out[5] sg13g2_tielo
XFILLER_25_217 VPWR VGND sg13g2_fill_2
XFILLER_33_250 VPWR VGND sg13g2_fill_2
X_4825_ _1749_ _1769_ _1771_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_957 VPWR VGND sg13g2_decap_8
X_4756_ _1701_ _1691_ _1703_ VPWR VGND sg13g2_xor2_1
X_3707_ _0867_ _0865_ _0866_ VPWR VGND sg13g2_nand2_1
X_4687_ _1634_ _1627_ _1635_ VPWR VGND sg13g2_xor2_1
X_3638_ net574 _0802_ _0803_ _0804_ _0805_ VPWR VGND sg13g2_nor4_1
X_3569_ VPWR VGND _0622_ _0736_ _0739_ net571 _0740_ _0701_ sg13g2_a221oi_1
X_5308_ net85 VGND VPWR _0067_ ppwm_i.u_ppwm.pc\[1\] clknet_leaf_21_clk sg13g2_dfrbpq_2
X_5239_ _2144_ falu_i.falutop.data_in\[14\] _2145_ VPWR VGND sg13g2_xor2_1
XFILLER_29_512 VPWR VGND sg13g2_decap_4
XFILLER_17_43 VPWR VGND sg13g2_decap_4
XFILLER_40_710 VPWR VGND sg13g2_decap_8
XFILLER_13_957 VPWR VGND sg13g2_decap_8
XFILLER_3_198 VPWR VGND sg13g2_fill_2
XFILLER_0_883 VPWR VGND sg13g2_decap_8
Xhold5 _0065_ VPWR VGND net377 sg13g2_dlygate4sd3_1
XFILLER_48_865 VPWR VGND sg13g2_decap_8
XFILLER_16_751 VPWR VGND sg13g2_fill_1
X_5290__117 VPWR VGND net117 sg13g2_tiehi
X_2940_ _2294_ net806 VPWR VGND sg13g2_inv_2
XFILLER_31_721 VPWR VGND sg13g2_decap_4
X_2871_ _2225_ net928 VPWR VGND sg13g2_inv_2
X_4610_ _1559_ _1553_ _1557_ _1558_ VPWR VGND sg13g2_and3_1
XFILLER_8_972 VPWR VGND sg13g2_decap_8
X_4541_ VGND VPWR _1487_ _1488_ _1491_ _1429_ sg13g2_a21oi_1
Xhold416 _0040_ VPWR VGND net1068 sg13g2_dlygate4sd3_1
XFILLER_7_493 VPWR VGND sg13g2_fill_2
Xhold427 falu_i.falutop.div_inst.rem\[7\] VPWR VGND net1079 sg13g2_dlygate4sd3_1
Xhold405 falu_i.falutop.i2c_inst.result\[1\] VPWR VGND net1057 sg13g2_dlygate4sd3_1
X_4472_ _1423_ _1397_ _1422_ VPWR VGND sg13g2_nand2_1
X_3423_ _0589_ VPWR _0601_ VGND _0599_ _0600_ sg13g2_o21ai_1
Xhold438 ppwm_i.u_ppwm.u_pwm.counter\[4\] VPWR VGND net1090 sg13g2_dlygate4sd3_1
Xhold449 falu_i.falutop.data_in\[11\] VPWR VGND net1101 sg13g2_dlygate4sd3_1
X_3354_ net581 _0531_ _0529_ _0532_ VPWR VGND sg13g2_nand3_1
XFILLER_31_0 VPWR VGND sg13g2_decap_8
X_3285_ _0468_ ppwm_i.u_ppwm.u_pwm.cmp_value\[5\] _2276_ ppwm_i.u_ppwm.u_pwm.cmp_value\[6\]
+ _2275_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_331 VPWR VGND sg13g2_decap_8
X_5024_ _1965_ VPWR _1966_ VGND _1919_ _1921_ sg13g2_o21ai_1
XFILLER_16_1007 VPWR VGND sg13g2_decap_8
XFILLER_21_242 VPWR VGND sg13g2_fill_1
X_4808_ _1754_ _1688_ _1751_ VPWR VGND sg13g2_nand2_1
X_4739_ _1633_ VPWR _1686_ VGND _1627_ _1634_ sg13g2_o21ai_1
XFILLER_1_603 VPWR VGND sg13g2_fill_1
XFILLER_1_658 VPWR VGND sg13g2_fill_1
X_5314__73 VPWR VGND net73 sg13g2_tiehi
XFILLER_49_618 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_fill_1
X_5360__332 VPWR VGND net332 sg13g2_tiehi
XFILLER_44_63 VPWR VGND sg13g2_fill_2
XFILLER_13_743 VPWR VGND sg13g2_fill_2
XFILLER_40_562 VPWR VGND sg13g2_fill_1
XFILLER_40_551 VPWR VGND sg13g2_fill_2
XFILLER_13_765 VPWR VGND sg13g2_decap_4
XFILLER_5_35 VPWR VGND sg13g2_fill_2
XFILLER_5_986 VPWR VGND sg13g2_decap_8
X_5406__240 VPWR VGND net240 sg13g2_tiehi
X_3070_ _2424_ _2423_ _2308_ VPWR VGND sg13g2_nand2b_1
XFILLER_36_857 VPWR VGND sg13g2_decap_4
X_3972_ VGND VPWR _2160_ net673 _0205_ _1014_ sg13g2_a21oi_1
X_2923_ VPWR _2277_ net1090 VGND sg13g2_inv_1
X_2854_ VPWR _2208_ net422 VGND sg13g2_inv_1
X_5573_ net40 VGND VPWR net968 falu_i.falutop.div_inst.b\[3\] clknet_leaf_3_clk sg13g2_dfrbpq_1
Xhold202 ppwm_i.u_ppwm.u_mem.memory\[43\] VPWR VGND net854 sg13g2_dlygate4sd3_1
X_4524_ _1473_ _1464_ _1474_ VPWR VGND sg13g2_xor2_1
Xhold235 falu_i.falutop.div_inst.start VPWR VGND net887 sg13g2_dlygate4sd3_1
Xhold224 _0119_ VPWR VGND net876 sg13g2_dlygate4sd3_1
Xhold213 _0044_ VPWR VGND net865 sg13g2_dlygate4sd3_1
X_4455_ _1407_ net939 _1405_ VPWR VGND sg13g2_xnor2_1
Xhold257 _0243_ VPWR VGND net909 sg13g2_dlygate4sd3_1
Xhold268 falu_i.falutop.div_inst.b\[6\] VPWR VGND net920 sg13g2_dlygate4sd3_1
Xhold246 ppwm_i.u_ppwm.u_mem.memory\[18\] VPWR VGND net898 sg13g2_dlygate4sd3_1
X_3406_ _0581_ _0582_ _0580_ _0584_ VPWR VGND _0583_ sg13g2_nand4_1
Xfanout704 _2306_ net704 VPWR VGND sg13g2_buf_8
Xhold279 falu_i.falutop.div_inst.acc\[6\] VPWR VGND net931 sg13g2_dlygate4sd3_1
Xfanout715 falu_i.falutop.alu_data_in\[15\] net715 VPWR VGND sg13g2_buf_8
X_4386_ VGND VPWR net743 net707 _1339_ net735 sg13g2_a21oi_1
X_3337_ VPWR _0069_ _0515_ VGND sg13g2_inv_1
Xfanout748 net749 net748 VPWR VGND sg13g2_buf_8
Xfanout726 falu_i.falutop.alu_data_in\[12\] net726 VPWR VGND sg13g2_buf_8
Xfanout737 net738 net737 VPWR VGND sg13g2_buf_8
Xfanout759 net760 net759 VPWR VGND sg13g2_buf_1
X_3268_ VGND VPWR ppwm_i.u_ppwm.global_counter\[16\] _0452_ _0454_ net989 sg13g2_a21oi_1
X_5457__58 VPWR VGND net58 sg13g2_tiehi
X_3199_ VGND VPWR _0409_ _0407_ _2277_ sg13g2_or2_1
X_5007_ net711 VPWR _1949_ VGND net768 net752 sg13g2_o21ai_1
XFILLER_38_183 VPWR VGND sg13g2_fill_1
XFILLER_26_323 VPWR VGND sg13g2_fill_2
XFILLER_26_378 VPWR VGND sg13g2_fill_2
XFILLER_14_66 VPWR VGND sg13g2_fill_1
X_5388__276 VPWR VGND net276 sg13g2_tiehi
XFILLER_2_967 VPWR VGND sg13g2_decap_8
XFILLER_49_448 VPWR VGND sg13g2_decap_8
XFILLER_18_802 VPWR VGND sg13g2_fill_1
XFILLER_18_879 VPWR VGND sg13g2_decap_8
XFILLER_29_194 VPWR VGND sg13g2_fill_2
XFILLER_45_676 VPWR VGND sg13g2_decap_4
XFILLER_44_197 VPWR VGND sg13g2_decap_8
XFILLER_13_540 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_13_595 VPWR VGND sg13g2_fill_1
XFILLER_9_588 VPWR VGND sg13g2_fill_2
XFILLER_9_599 VPWR VGND sg13g2_fill_2
X_4240_ VGND VPWR net605 _1201_ _0285_ _1202_ sg13g2_a21oi_1
X_4171_ VGND VPWR _2149_ net636 _0268_ _1150_ sg13g2_a21oi_1
X_3122_ VGND VPWR net802 _0357_ _0011_ _0358_ sg13g2_a21oi_1
XFILLER_49_971 VPWR VGND sg13g2_decap_8
X_3053_ VPWR VGND _2163_ _2405_ net695 _2158_ _2407_ net702 sg13g2_a221oi_1
XFILLER_24_816 VPWR VGND sg13g2_decap_8
XFILLER_17_890 VPWR VGND sg13g2_decap_8
X_3955_ net841 VPWR _1006_ VGND net961 net674 sg13g2_o21ai_1
X_2906_ VPWR _2260_ ppwm_i.u_ppwm.global_counter\[17\] VGND sg13g2_inv_1
X_3886_ VGND VPWR _2191_ net670 _0162_ _0971_ sg13g2_a21oi_1
X_2837_ VPWR _2191_ net491 VGND sg13g2_inv_1
X_5556_ net210 VGND VPWR net1128 falu_i.falutop.alu_data_in\[2\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_4507_ _1404_ VPWR _1458_ VGND net939 falu_i.falutop.div_inst.val\[0\] sg13g2_o21ai_1
X_5487_ net309 VGND VPWR _0246_ falu_i.falutop.div_inst.quo\[0\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_5528__161 VPWR VGND net161 sg13g2_tiehi
X_4438_ _1387_ _1388_ _1382_ _1390_ VPWR VGND _1389_ sg13g2_nand4_1
X_4369_ _1260_ _1321_ _1322_ VPWR VGND sg13g2_nor2_2
XFILLER_46_407 VPWR VGND sg13g2_fill_1
Xfanout578 net580 net578 VPWR VGND sg13g2_buf_1
Xfanout589 net590 net589 VPWR VGND sg13g2_buf_8
Xfanout567 net568 net567 VPWR VGND sg13g2_buf_8
XFILLER_30_808 VPWR VGND sg13g2_fill_1
XFILLER_41_20 VPWR VGND sg13g2_fill_1
XFILLER_10_554 VPWR VGND sg13g2_decap_4
XFILLER_10_587 VPWR VGND sg13g2_fill_2
XFILLER_6_569 VPWR VGND sg13g2_decap_4
XFILLER_2_720 VPWR VGND sg13g2_fill_2
XFILLER_29_1028 VPWR VGND sg13g2_fill_1
XFILLER_46_930 VPWR VGND sg13g2_decap_8
XFILLER_18_632 VPWR VGND sg13g2_fill_2
XFILLER_45_473 VPWR VGND sg13g2_decap_8
XFILLER_17_164 VPWR VGND sg13g2_fill_2
XFILLER_21_819 VPWR VGND sg13g2_decap_8
X_3740_ _0895_ _0896_ net575 _0897_ VPWR VGND sg13g2_nand3_1
XFILLER_20_307 VPWR VGND sg13g2_fill_1
XFILLER_12_1021 VPWR VGND sg13g2_decap_8
X_3671_ net577 VPWR _0835_ VGND ppwm_i.u_ppwm.pwm_value\[2\] net582 sg13g2_o21ai_1
X_5410_ net232 VGND VPWR net464 ppwm_i.u_ppwm.u_mem.memory\[69\] clknet_leaf_27_clk
+ sg13g2_dfrbpq_1
X_5341_ net370 VGND VPWR _0100_ ppwm_i.u_ppwm.u_mem.memory\[0\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
X_5272_ net152 VGND VPWR net1113 ppwm_i.u_ppwm.u_pwm.counter\[0\] clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
X_4223_ net411 net605 _1190_ VPWR VGND sg13g2_nor2_1
X_4154_ _1144_ _1104_ net994 net967 net778 VPWR VGND sg13g2_a22oi_1
X_4085_ _1089_ _2438_ falu_i.falutop.i2c_inst.result\[4\] _2432_ falu_i.falutop.i2c_inst.result\[7\]
+ VPWR VGND sg13g2_a22oi_1
X_3105_ VGND VPWR net801 _0345_ _0006_ _0346_ sg13g2_a21oi_1
X_3036_ VGND VPWR _2390_ net612 net603 sg13g2_or2_1
XFILLER_37_985 VPWR VGND sg13g2_decap_8
XFILLER_24_624 VPWR VGND sg13g2_decap_8
XFILLER_36_484 VPWR VGND sg13g2_fill_1
XFILLER_23_134 VPWR VGND sg13g2_decap_8
XFILLER_24_657 VPWR VGND sg13g2_decap_8
X_4987_ _1930_ falu_i.falutop.div_inst.rem\[2\] _1928_ VPWR VGND sg13g2_xnor2_1
XFILLER_23_189 VPWR VGND sg13g2_fill_1
X_5450__86 VPWR VGND net86 sg13g2_tiehi
X_3938_ VGND VPWR _2172_ net667 _0188_ _0997_ sg13g2_a21oi_1
X_3869_ net825 VPWR _0963_ VGND net398 net645 sg13g2_o21ai_1
XFILLER_20_874 VPWR VGND sg13g2_decap_8
XFILLER_3_517 VPWR VGND sg13g2_decap_4
X_5539_ net68 VGND VPWR _0298_ falu_i.falutop.i2c_inst.result\[3\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
XFILLER_28_952 VPWR VGND sg13g2_decap_8
XFILLER_43_933 VPWR VGND sg13g2_decap_8
XFILLER_15_613 VPWR VGND sg13g2_fill_1
XFILLER_27_473 VPWR VGND sg13g2_fill_1
XFILLER_14_167 VPWR VGND sg13g2_decap_8
XFILLER_6_311 VPWR VGND sg13g2_decap_8
XFILLER_11_874 VPWR VGND sg13g2_decap_8
XFILLER_7_867 VPWR VGND sg13g2_decap_8
XFILLER_6_322 VPWR VGND sg13g2_fill_2
XFILLER_6_399 VPWR VGND sg13g2_fill_2
XFILLER_2_550 VPWR VGND sg13g2_fill_2
X_4910_ _1854_ net723 _1803_ VPWR VGND sg13g2_nand2_1
XFILLER_19_996 VPWR VGND sg13g2_decap_8
XFILLER_45_292 VPWR VGND sg13g2_fill_2
X_4841_ _1723_ VPWR _1786_ VGND net705 _1654_ sg13g2_o21ai_1
XFILLER_34_955 VPWR VGND sg13g2_decap_8
X_4772_ _1650_ _1718_ _0301_ VPWR VGND sg13g2_nor2_1
X_3723_ VPWR VGND _0881_ net798 _0878_ _2236_ _0089_ net569 sg13g2_a221oi_1
X_3654_ _0813_ _0819_ _0636_ _0820_ VPWR VGND sg13g2_nand3_1
X_3585_ net574 _0753_ _0754_ _0755_ VPWR VGND sg13g2_nor3_1
X_5324_ net53 VGND VPWR _0083_ ppwm_i.u_ppwm.u_ex.reg_value_q\[1\] clknet_leaf_8_clk
+ sg13g2_dfrbpq_2
X_5255_ net185 VGND VPWR _0017_ falu_i.falutop.i2c_inst.data_in\[13\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_4206_ VGND VPWR net633 _1175_ _0277_ _1176_ sg13g2_a21oi_1
X_5186_ net1086 net617 _2108_ VPWR VGND sg13g2_nor2_1
X_4137_ _0248_ _2298_ net619 net833 _2291_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_771 VPWR VGND sg13g2_decap_4
X_4068_ net899 falu_i.falutop.data_in\[9\] net685 _0237_ VPWR VGND sg13g2_mux2_1
XFILLER_25_911 VPWR VGND sg13g2_decap_8
XFILLER_37_782 VPWR VGND sg13g2_fill_1
X_3019_ VPWR VGND _2372_ net786 _2371_ _2368_ _2373_ _2369_ sg13g2_a221oi_1
XFILLER_40_925 VPWR VGND sg13g2_decap_8
XFILLER_40_914 VPWR VGND sg13g2_decap_8
XFILLER_25_988 VPWR VGND sg13g2_decap_8
XFILLER_11_126 VPWR VGND sg13g2_fill_2
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_20_682 VPWR VGND sg13g2_decap_4
XFILLER_22_99 VPWR VGND sg13g2_fill_1
XFILLER_4_859 VPWR VGND sg13g2_decap_8
XFILLER_16_944 VPWR VGND sg13g2_decap_8
XFILLER_15_432 VPWR VGND sg13g2_decap_8
XFILLER_15_443 VPWR VGND sg13g2_fill_1
X_5370__312 VPWR VGND net312 sg13g2_tiehi
XFILLER_31_947 VPWR VGND sg13g2_decap_8
XFILLER_7_620 VPWR VGND sg13g2_decap_8
XFILLER_11_671 VPWR VGND sg13g2_fill_1
X_3370_ _2243_ net596 _0548_ VPWR VGND sg13g2_nor2_1
X_5040_ _1878_ VPWR _1981_ VGND _1827_ _1877_ sg13g2_o21ai_1
Xheichips25_tiny_wrapper_28 VPWR VGND uo_out[6] sg13g2_tielo
Xheichips25_tiny_wrapper_17 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_19_782 VPWR VGND sg13g2_fill_1
XFILLER_46_590 VPWR VGND sg13g2_fill_1
XFILLER_34_752 VPWR VGND sg13g2_fill_2
X_5416__220 VPWR VGND net220 sg13g2_tiehi
XFILLER_22_936 VPWR VGND sg13g2_decap_8
XFILLER_33_262 VPWR VGND sg13g2_fill_2
X_4824_ _1770_ _1749_ _1769_ VPWR VGND sg13g2_nand2b_1
X_4755_ _1699_ _1700_ _1691_ _1702_ VPWR VGND sg13g2_nand3_1
X_3706_ _0866_ _0850_ _0856_ VPWR VGND sg13g2_nand2_1
X_4686_ _1632_ _1628_ _1634_ VPWR VGND sg13g2_xor2_1
X_3637_ _0701_ _0714_ _0804_ VPWR VGND sg13g2_nor2_1
X_3568_ VGND VPWR net610 _0738_ _0739_ _0737_ sg13g2_a21oi_1
X_5307_ net87 VGND VPWR net1164 ppwm_i.u_ppwm.pc\[0\] clknet_leaf_23_clk sg13g2_dfrbpq_2
X_5347__358 VPWR VGND net358 sg13g2_tiehi
X_3499_ _0673_ net611 _0651_ VPWR VGND sg13g2_nand2_1
X_5238_ _2144_ net773 _2093_ VPWR VGND sg13g2_nand2_1
X_5169_ net1141 net620 _2103_ VPWR VGND sg13g2_nor2_1
XFILLER_17_719 VPWR VGND sg13g2_fill_2
XFILLER_13_936 VPWR VGND sg13g2_decap_8
XFILLER_24_273 VPWR VGND sg13g2_fill_2
XFILLER_33_32 VPWR VGND sg13g2_fill_1
XFILLER_12_457 VPWR VGND sg13g2_fill_1
XFILLER_21_980 VPWR VGND sg13g2_decap_8
XFILLER_32_1024 VPWR VGND sg13g2_decap_4
XFILLER_4_634 VPWR VGND sg13g2_decap_8
XFILLER_4_623 VPWR VGND sg13g2_fill_1
XFILLER_4_612 VPWR VGND sg13g2_decap_8
XFILLER_4_656 VPWR VGND sg13g2_fill_1
XFILLER_4_689 VPWR VGND sg13g2_fill_2
XFILLER_0_862 VPWR VGND sg13g2_decap_8
Xhold6 ppwm_i.u_ppwm.u_mem.bit_count\[0\] VPWR VGND net378 sg13g2_dlygate4sd3_1
XFILLER_47_332 VPWR VGND sg13g2_fill_1
X_5398__256 VPWR VGND net256 sg13g2_tiehi
XFILLER_16_730 VPWR VGND sg13g2_fill_2
XFILLER_15_240 VPWR VGND sg13g2_fill_1
X_2870_ VPWR _2224_ net496 VGND sg13g2_inv_1
XFILLER_8_951 VPWR VGND sg13g2_decap_8
X_4540_ _1487_ _1488_ _1429_ _1490_ VPWR VGND sg13g2_nand3_1
Xclkbuf_leaf_10_clk clknet_3_3__leaf_clk clknet_leaf_10_clk VPWR VGND sg13g2_buf_8
Xhold406 _0296_ VPWR VGND net1058 sg13g2_dlygate4sd3_1
X_4471_ _1422_ _1414_ _1420_ VPWR VGND sg13g2_xnor2_1
Xhold417 falu_i.falutop.i2c_inst.data_in\[19\] VPWR VGND net1069 sg13g2_dlygate4sd3_1
X_3422_ _2243_ ppwm_i.u_ppwm.global_counter\[19\] _0600_ VPWR VGND sg13g2_nor2_1
Xhold439 _0038_ VPWR VGND net1091 sg13g2_dlygate4sd3_1
Xhold428 _1184_ VPWR VGND net1080 sg13g2_dlygate4sd3_1
X_3353_ VGND VPWR _2235_ ppwm_i.u_ppwm.pwm_value\[9\] _0531_ net591 sg13g2_a21oi_1
X_3284_ _2283_ ppwm_i.u_ppwm.u_pwm.counter\[5\] _0466_ _0467_ VPWR VGND sg13g2_a21o_1
XFILLER_24_0 VPWR VGND sg13g2_fill_2
X_5023_ VPWR _1965_ _1964_ VGND sg13g2_inv_1
XFILLER_26_505 VPWR VGND sg13g2_fill_1
XFILLER_19_590 VPWR VGND sg13g2_decap_8
X_4807_ _1753_ net713 net768 VPWR VGND sg13g2_nand2_1
X_2999_ VGND VPWR _2351_ _2352_ _2353_ _2254_ sg13g2_a21oi_1
XFILLER_21_276 VPWR VGND sg13g2_fill_1
X_4738_ _1683_ _1682_ _1685_ VPWR VGND sg13g2_xor2_1
X_4669_ _1615_ _1616_ _1614_ _1617_ VPWR VGND sg13g2_nand3_1
XFILLER_28_21 VPWR VGND sg13g2_decap_8
XFILLER_17_516 VPWR VGND sg13g2_decap_8
XFILLER_17_527 VPWR VGND sg13g2_fill_2
XFILLER_12_243 VPWR VGND sg13g2_decap_8
XFILLER_9_748 VPWR VGND sg13g2_decap_4
XFILLER_8_247 VPWR VGND sg13g2_decap_4
XFILLER_5_965 VPWR VGND sg13g2_decap_8
XFILLER_4_464 VPWR VGND sg13g2_fill_2
XFILLER_0_681 VPWR VGND sg13g2_fill_1
XFILLER_0_692 VPWR VGND sg13g2_decap_8
XFILLER_39_1008 VPWR VGND sg13g2_decap_8
XFILLER_16_560 VPWR VGND sg13g2_fill_1
X_3971_ net837 VPWR _1014_ VGND ppwm_i.u_ppwm.u_mem.memory\[105\] net673 sg13g2_o21ai_1
X_2922_ VPWR _2276_ net1060 VGND sg13g2_inv_1
X_2853_ VPWR _2207_ net455 VGND sg13g2_inv_1
X_5572_ net48 VGND VPWR net892 falu_i.falutop.div_inst.b\[2\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_8_781 VPWR VGND sg13g2_decap_8
XFILLER_8_770 VPWR VGND sg13g2_decap_8
X_4523_ _1473_ _1465_ _1471_ VPWR VGND sg13g2_xnor2_1
Xhold203 _0142_ VPWR VGND net855 sg13g2_dlygate4sd3_1
Xhold214 ppwm_i.u_ppwm.u_mem.memory\[59\] VPWR VGND net866 sg13g2_dlygate4sd3_1
Xhold225 falu_i.falutop.alu_inst.op\[0\] VPWR VGND net877 sg13g2_dlygate4sd3_1
X_4454_ _1406_ net380 net639 VPWR VGND sg13g2_nand2_2
Xhold258 falu_i.falutop.div_inst.quo\[0\] VPWR VGND net910 sg13g2_dlygate4sd3_1
Xhold269 _0335_ VPWR VGND net921 sg13g2_dlygate4sd3_1
Xhold247 falu_i.falutop.i2c_inst.data_in\[9\] VPWR VGND net899 sg13g2_dlygate4sd3_1
Xhold236 ppwm_i.u_ppwm.u_mem.memory\[11\] VPWR VGND net888 sg13g2_dlygate4sd3_1
X_3405_ _0583_ _2260_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] _2259_ net782 VPWR VGND
+ sg13g2_a22oi_1
X_5266__164 VPWR VGND net164 sg13g2_tiehi
Xfanout705 _2302_ net705 VPWR VGND sg13g2_buf_8
X_4385_ VPWR _1338_ _1337_ VGND sg13g2_inv_1
X_3336_ _0515_ _0513_ _0514_ _0493_ net786 VPWR VGND sg13g2_a22oi_1
Xfanout716 net717 net716 VPWR VGND sg13g2_buf_8
Xfanout738 net739 net738 VPWR VGND sg13g2_buf_8
Xfanout727 net729 net727 VPWR VGND sg13g2_buf_8
Xfanout749 net1131 net749 VPWR VGND sg13g2_buf_8
X_3267_ net796 net1126 _0061_ VPWR VGND sg13g2_nor2_1
X_5006_ VPWR _1948_ _1947_ VGND sg13g2_inv_1
X_3198_ VGND VPWR _2278_ net1050 _0037_ _0408_ sg13g2_a21oi_1
XFILLER_38_195 VPWR VGND sg13g2_decap_4
XFILLER_14_78 VPWR VGND sg13g2_fill_1
XFILLER_2_946 VPWR VGND sg13g2_decap_8
XFILLER_49_405 VPWR VGND sg13g2_decap_8
XFILLER_49_427 VPWR VGND sg13g2_decap_8
XFILLER_7_1028 VPWR VGND sg13g2_fill_1
X_5579__263 VPWR VGND net263 sg13g2_tiehi
XFILLER_18_858 VPWR VGND sg13g2_decap_8
XFILLER_44_143 VPWR VGND sg13g2_fill_1
XFILLER_32_305 VPWR VGND sg13g2_fill_2
XFILLER_44_187 VPWR VGND sg13g2_fill_1
XFILLER_13_574 VPWR VGND sg13g2_decap_8
XFILLER_5_773 VPWR VGND sg13g2_fill_2
X_4170_ net818 VPWR _1150_ VGND net905 net636 sg13g2_o21ai_1
X_3121_ net804 VPWR _0358_ VGND net871 _0357_ sg13g2_o21ai_1
XFILLER_49_950 VPWR VGND sg13g2_decap_8
X_3052_ VGND VPWR _2168_ net690 _2406_ net709 sg13g2_a21oi_1
XFILLER_35_154 VPWR VGND sg13g2_fill_1
XFILLER_35_198 VPWR VGND sg13g2_decap_8
X_3954_ VGND VPWR _2167_ net649 _0196_ _1005_ sg13g2_a21oi_1
XFILLER_16_390 VPWR VGND sg13g2_fill_1
X_2905_ _2259_ net1076 VPWR VGND sg13g2_inv_2
X_3885_ net834 VPWR _0971_ VGND net474 net670 sg13g2_o21ai_1
XFILLER_32_883 VPWR VGND sg13g2_fill_2
X_2836_ VPWR _2190_ net449 VGND sg13g2_inv_1
X_5555_ net215 VGND VPWR net1142 falu_i.falutop.alu_data_in\[1\] clknet_leaf_35_clk
+ sg13g2_dfrbpq_1
X_5486_ net311 VGND VPWR _0245_ falu_i.falutop.div_inst.acc\[0\] clknet_leaf_44_clk
+ sg13g2_dfrbpq_2
X_4506_ net818 VPWR _1457_ VGND net1047 net628 sg13g2_o21ai_1
XFILLER_6_90 VPWR VGND sg13g2_decap_8
X_4437_ VGND VPWR _1232_ _1319_ _1389_ _1381_ sg13g2_a21oi_1
X_4368_ _1321_ falu_i.falutop.alu_inst.op\[2\] _2300_ VPWR VGND sg13g2_nand2_2
Xfanout579 net580 net579 VPWR VGND sg13g2_buf_8
X_3319_ _0499_ _0496_ _0498_ VPWR VGND sg13g2_xnor2_1
Xfanout568 _1132_ net568 VPWR VGND sg13g2_buf_8
X_4299_ _1252_ _1235_ _1250_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_338 VPWR VGND sg13g2_decap_8
XFILLER_25_44 VPWR VGND sg13g2_decap_4
XFILLER_41_146 VPWR VGND sg13g2_decap_8
XFILLER_41_179 VPWR VGND sg13g2_decap_8
XFILLER_10_533 VPWR VGND sg13g2_decap_4
XFILLER_41_65 VPWR VGND sg13g2_fill_2
XFILLER_41_43 VPWR VGND sg13g2_fill_2
XFILLER_2_710 VPWR VGND sg13g2_fill_2
X_5507__257 VPWR VGND net257 sg13g2_tiehi
XFILLER_2_765 VPWR VGND sg13g2_fill_1
XFILLER_2_787 VPWR VGND sg13g2_decap_8
XFILLER_37_408 VPWR VGND sg13g2_fill_1
XFILLER_46_986 VPWR VGND sg13g2_decap_8
XFILLER_17_143 VPWR VGND sg13g2_fill_1
XFILLER_18_688 VPWR VGND sg13g2_decap_8
XFILLER_14_894 VPWR VGND sg13g2_decap_8
XFILLER_9_353 VPWR VGND sg13g2_fill_2
XFILLER_12_1000 VPWR VGND sg13g2_decap_8
X_3670_ _0834_ net576 _0832_ _0833_ VPWR VGND sg13g2_and3_1
X_5340_ net371 VGND VPWR _0099_ ppwm_i.u_ppwm.u_mem.data_sync1 clknet_leaf_11_clk
+ sg13g2_dfrbpq_1
X_5271_ net154 VGND VPWR net536 ppwm_i.u_ppwm.u_pwm.cmp_value\[9\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
X_4222_ VGND VPWR net780 net388 _1189_ _1188_ sg13g2_a21oi_1
X_4153_ net1059 net891 _1103_ _0257_ VPWR VGND sg13g2_mux2_1
X_4084_ _1088_ _2430_ _1087_ VPWR VGND sg13g2_nand2_1
X_3104_ net820 VPWR _0346_ VGND net972 _0345_ sg13g2_o21ai_1
X_3035_ _2381_ _2388_ _2389_ VPWR VGND sg13g2_nor2_1
XFILLER_37_964 VPWR VGND sg13g2_decap_8
XFILLER_36_430 VPWR VGND sg13g2_fill_1
XFILLER_36_474 VPWR VGND sg13g2_fill_1
X_4986_ _1929_ _1928_ falu_i.falutop.div_inst.rem\[2\] VPWR VGND sg13g2_nand2b_1
X_3937_ net836 VPWR _0997_ VGND net541 net668 sg13g2_o21ai_1
X_3868_ VGND VPWR _2197_ net657 _0153_ _0962_ sg13g2_a21oi_1
XFILLER_20_853 VPWR VGND sg13g2_decap_8
X_3799_ net824 VPWR _0928_ VGND ppwm_i.u_ppwm.u_mem.memory\[20\] net641 sg13g2_o21ai_1
X_2819_ VPWR _2173_ net518 VGND sg13g2_inv_1
XFILLER_11_46 VPWR VGND sg13g2_fill_2
X_5538_ net76 VGND VPWR net1048 falu_i.falutop.i2c_inst.result\[2\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_5469_ net347 VGND VPWR net849 falu_i.falutop.data_in\[0\] clknet_leaf_8_clk sg13g2_dfrbpq_2
XFILLER_47_706 VPWR VGND sg13g2_fill_1
XFILLER_28_931 VPWR VGND sg13g2_decap_8
XFILLER_27_463 VPWR VGND sg13g2_fill_1
XFILLER_15_625 VPWR VGND sg13g2_fill_2
X_5357__338 VPWR VGND net338 sg13g2_tiehi
XFILLER_42_455 VPWR VGND sg13g2_fill_2
XFILLER_43_989 VPWR VGND sg13g2_decap_8
XFILLER_42_488 VPWR VGND sg13g2_fill_1
XFILLER_11_853 VPWR VGND sg13g2_decap_8
XFILLER_7_846 VPWR VGND sg13g2_decap_8
XFILLER_6_356 VPWR VGND sg13g2_fill_1
XFILLER_42_1015 VPWR VGND sg13g2_decap_8
XFILLER_38_706 VPWR VGND sg13g2_fill_1
XFILLER_37_238 VPWR VGND sg13g2_decap_4
XFILLER_19_975 VPWR VGND sg13g2_decap_8
XFILLER_34_934 VPWR VGND sg13g2_decap_8
X_4840_ _1784_ _1785_ _0302_ VPWR VGND sg13g2_nor2_1
X_4771_ VPWR VGND net639 net630 _1717_ net614 _1718_ _1715_ sg13g2_a221oi_1
X_3722_ _0774_ net569 _0880_ _0881_ VPWR VGND sg13g2_nor3_1
XFILLER_13_190 VPWR VGND sg13g2_fill_1
XFILLER_20_149 VPWR VGND sg13g2_fill_1
X_3653_ VPWR VGND net576 _0638_ _0818_ net579 _0819_ _0817_ sg13g2_a221oi_1
X_3584_ net584 _0647_ _0754_ VPWR VGND sg13g2_nor2_1
X_5323_ net55 VGND VPWR _0082_ ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_2
X_5254_ net187 VGND VPWR _0016_ falu_i.falutop.i2c_inst.data_in\[12\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_4205_ net803 VPWR _1176_ VGND net1106 net634 sg13g2_o21ai_1
X_5185_ net1103 net725 net617 _0325_ VPWR VGND sg13g2_mux2_1
X_4136_ _1136_ net820 _1074_ VPWR VGND sg13g2_nand2_1
XFILLER_29_717 VPWR VGND sg13g2_decap_4
X_4067_ net873 falu_i.falutop.data_in\[8\] net684 _0236_ VPWR VGND sg13g2_mux2_1
X_3018_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[34\] _2370_ net696 ppwm_i.u_ppwm.u_mem.memory\[55\]
+ _2372_ net700 sg13g2_a221oi_1
XFILLER_19_1017 VPWR VGND sg13g2_decap_8
XFILLER_25_967 VPWR VGND sg13g2_decap_8
XFILLER_19_1028 VPWR VGND sg13g2_fill_1
XFILLER_24_466 VPWR VGND sg13g2_fill_2
X_4969_ _1911_ _1906_ _1912_ VPWR VGND sg13g2_xor2_1
XFILLER_22_67 VPWR VGND sg13g2_fill_2
XFILLER_22_78 VPWR VGND sg13g2_fill_2
XFILLER_4_838 VPWR VGND sg13g2_decap_8
XFILLER_28_761 VPWR VGND sg13g2_fill_1
XFILLER_16_923 VPWR VGND sg13g2_decap_8
X_5474__337 VPWR VGND net337 sg13g2_tiehi
XFILLER_42_274 VPWR VGND sg13g2_fill_2
XFILLER_8_36 VPWR VGND sg13g2_fill_1
X_5568__80 VPWR VGND net80 sg13g2_tiehi
XFILLER_30_469 VPWR VGND sg13g2_decap_8
XFILLER_3_882 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_4
Xheichips25_tiny_wrapper_29 VPWR VGND uo_out[7] sg13g2_tielo
Xheichips25_tiny_wrapper_18 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_34_720 VPWR VGND sg13g2_fill_2
XFILLER_46_580 VPWR VGND sg13g2_decap_4
XFILLER_18_271 VPWR VGND sg13g2_fill_2
XFILLER_22_915 VPWR VGND sg13g2_decap_8
XFILLER_33_252 VPWR VGND sg13g2_fill_1
X_4823_ _1769_ _1757_ _1768_ VPWR VGND sg13g2_xnor2_1
X_4754_ _1701_ _1699_ _1700_ VPWR VGND sg13g2_nand2_1
X_3705_ net600 VPWR _0865_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[5\] ppwm_i.u_ppwm.u_ex.reg_value_q\[4\]
+ sg13g2_o21ai_1
X_4685_ _1633_ _1628_ _1632_ VPWR VGND sg13g2_nand2b_1
X_3636_ _0647_ _0694_ _0803_ VPWR VGND sg13g2_nor2_1
X_3567_ VGND VPWR ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] net596 _0738_ _0548_ sg13g2_a21oi_1
XFILLER_1_819 VPWR VGND sg13g2_decap_8
X_5306_ net88 VGND VPWR net1040 ppwm_i.u_ppwm.u_ex.state_q\[2\] clknet_leaf_18_clk
+ sg13g2_dfrbpq_2
X_5237_ net439 net625 _2143_ VPWR VGND sg13g2_nor2_1
X_3498_ _0671_ VPWR _0672_ VGND _0668_ _0669_ sg13g2_o21ai_1
X_5168_ VGND VPWR _2301_ net620 _0313_ _2102_ sg13g2_a21oi_1
X_5099_ _2038_ _2037_ _2039_ VPWR VGND sg13g2_xor2_1
X_4119_ _1120_ _1119_ _1115_ _1121_ VPWR VGND sg13g2_a21o_1
XFILLER_17_709 VPWR VGND sg13g2_fill_1
XFILLER_29_558 VPWR VGND sg13g2_fill_2
XFILLER_44_517 VPWR VGND sg13g2_fill_1
X_5276__144 VPWR VGND net144 sg13g2_tiehi
XFILLER_25_742 VPWR VGND sg13g2_decap_8
XFILLER_13_915 VPWR VGND sg13g2_decap_8
XFILLER_24_252 VPWR VGND sg13g2_fill_2
XFILLER_25_786 VPWR VGND sg13g2_fill_1
XFILLER_40_756 VPWR VGND sg13g2_fill_2
XFILLER_32_1003 VPWR VGND sg13g2_decap_8
XFILLER_20_491 VPWR VGND sg13g2_decap_8
XFILLER_0_841 VPWR VGND sg13g2_decap_8
XFILLER_48_812 VPWR VGND sg13g2_fill_2
Xhold7 _0212_ VPWR VGND net379 sg13g2_dlygate4sd3_1
XFILLER_43_561 VPWR VGND sg13g2_fill_1
XFILLER_30_211 VPWR VGND sg13g2_fill_2
XFILLER_8_930 VPWR VGND sg13g2_decap_8
XFILLER_11_491 VPWR VGND sg13g2_decap_8
X_4470_ _1421_ _1420_ _1414_ VPWR VGND sg13g2_nand2b_1
Xhold407 falu_i.falutop.div_inst.b1\[2\] VPWR VGND net1059 sg13g2_dlygate4sd3_1
Xhold418 falu_i.falutop.i2c_inst.data_in\[16\] VPWR VGND net1070 sg13g2_dlygate4sd3_1
X_3421_ VGND VPWR _2244_ ppwm_i.u_ppwm.global_counter\[18\] _0599_ _0598_ sg13g2_a21oi_1
XFILLER_7_495 VPWR VGND sg13g2_fill_1
Xhold429 falu_i.falutop.div_inst.b\[0\] VPWR VGND net1081 sg13g2_dlygate4sd3_1
X_3352_ net612 _2419_ _0530_ VPWR VGND sg13g2_nor2_1
X_3283_ VGND VPWR _2277_ ppwm_i.u_ppwm.u_pwm.cmp_value\[4\] _0466_ _0465_ sg13g2_a21oi_1
X_5022_ _1964_ _1933_ _1962_ VPWR VGND sg13g2_xnor2_1
XFILLER_17_0 VPWR VGND sg13g2_decap_4
XFILLER_38_399 VPWR VGND sg13g2_fill_2
XFILLER_0_1023 VPWR VGND sg13g2_decap_4
XFILLER_22_745 VPWR VGND sg13g2_fill_2
X_4806_ _1752_ net711 net766 VPWR VGND sg13g2_nand2_2
XFILLER_10_929 VPWR VGND sg13g2_decap_8
XFILLER_22_789 VPWR VGND sg13g2_decap_8
X_2998_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[100\] net709 net694 ppwm_i.u_ppwm.u_mem.memory\[86\]
+ _2352_ net698 sg13g2_a221oi_1
X_4737_ _1684_ _1682_ _1683_ VPWR VGND sg13g2_nand2b_1
X_4668_ VGND VPWR _1218_ _1322_ _1616_ _1613_ sg13g2_a21oi_1
X_3619_ net585 _0700_ _0787_ VPWR VGND sg13g2_nor2_1
X_4599_ _1490_ VPWR _1548_ VGND _1482_ _1491_ sg13g2_o21ai_1
XFILLER_0_115 VPWR VGND sg13g2_decap_8
XFILLER_0_159 VPWR VGND sg13g2_decap_8
XFILLER_0_137 VPWR VGND sg13g2_fill_2
XFILLER_29_311 VPWR VGND sg13g2_decap_8
XFILLER_28_44 VPWR VGND sg13g2_fill_2
XFILLER_44_65 VPWR VGND sg13g2_fill_1
XFILLER_40_520 VPWR VGND sg13g2_fill_1
XFILLER_8_204 VPWR VGND sg13g2_decap_4
XFILLER_5_944 VPWR VGND sg13g2_decap_8
XFILLER_48_620 VPWR VGND sg13g2_decap_8
X_5521__190 VPWR VGND net190 sg13g2_tiehi
XFILLER_48_697 VPWR VGND sg13g2_fill_1
X_3970_ VGND VPWR _2161_ net673 _0204_ _1013_ sg13g2_a21oi_1
XFILLER_43_380 VPWR VGND sg13g2_decap_8
X_2921_ VPWR _2275_ net1066 VGND sg13g2_inv_1
X_2852_ VPWR _2206_ net969 VGND sg13g2_inv_1
X_5571_ net56 VGND VPWR net414 falu_i.falutop.div_inst.b\[1\] clknet_leaf_2_clk sg13g2_dfrbpq_1
X_4522_ _1472_ _1465_ _1471_ VPWR VGND sg13g2_nand2_1
Xhold215 ppwm_i.u_ppwm.u_mem.memory\[94\] VPWR VGND net867 sg13g2_dlygate4sd3_1
X_4453_ _1405_ falu_i.falutop.div_inst.val\[0\] _1404_ VPWR VGND sg13g2_nand2_1
Xhold204 falu_i.falutop.div_inst.acc\[4\] VPWR VGND net856 sg13g2_dlygate4sd3_1
Xhold226 ppwm_i.u_ppwm.u_mem.memory\[84\] VPWR VGND net878 sg13g2_dlygate4sd3_1
X_3404_ _0582_ ppwm_i.u_ppwm.global_counter\[18\] net782 VPWR VGND sg13g2_nand2b_1
Xhold237 ppwm_i.u_ppwm.u_mem.memory\[67\] VPWR VGND net889 sg13g2_dlygate4sd3_1
Xhold259 _1133_ VPWR VGND net911 sg13g2_dlygate4sd3_1
Xhold248 _0237_ VPWR VGND net900 sg13g2_dlygate4sd3_1
Xfanout706 _2302_ net706 VPWR VGND sg13g2_buf_1
X_4384_ net771 _1302_ _2299_ _1337_ VPWR VGND sg13g2_nand3_1
X_3335_ VPWR VGND _0482_ _2422_ _0510_ _0478_ _0514_ _0506_ sg13g2_a221oi_1
Xfanout717 net720 net717 VPWR VGND sg13g2_buf_8
Xfanout728 net729 net728 VPWR VGND sg13g2_buf_2
Xfanout739 falu_i.falutop.alu_data_in\[10\] net739 VPWR VGND sg13g2_buf_8
X_3266_ _0453_ net1125 _0452_ VPWR VGND sg13g2_xnor2_1
X_5005_ VGND VPWR _1944_ _1947_ _1907_ _1752_ sg13g2_a21oi_2
XFILLER_22_1013 VPWR VGND sg13g2_decap_8
XFILLER_39_664 VPWR VGND sg13g2_fill_2
X_3197_ _0408_ net809 _0407_ VPWR VGND sg13g2_nand2_1
XFILLER_14_509 VPWR VGND sg13g2_decap_8
XFILLER_14_57 VPWR VGND sg13g2_decap_8
XFILLER_22_575 VPWR VGND sg13g2_fill_1
XFILLER_10_737 VPWR VGND sg13g2_decap_8
XFILLER_10_748 VPWR VGND sg13g2_fill_1
XFILLER_2_925 VPWR VGND sg13g2_decap_8
X_5245__205 VPWR VGND net205 sg13g2_tiehi
XFILLER_7_1007 VPWR VGND sg13g2_decap_8
XFILLER_17_314 VPWR VGND sg13g2_decap_8
XFILLER_18_837 VPWR VGND sg13g2_decap_8
XFILLER_29_174 VPWR VGND sg13g2_fill_2
XFILLER_29_196 VPWR VGND sg13g2_fill_1
XFILLER_26_881 VPWR VGND sg13g2_decap_8
XFILLER_32_317 VPWR VGND sg13g2_fill_1
XFILLER_9_557 VPWR VGND sg13g2_decap_8
XFILLER_9_568 VPWR VGND sg13g2_fill_1
X_5367__318 VPWR VGND net318 sg13g2_tiehi
XFILLER_5_763 VPWR VGND sg13g2_fill_1
XFILLER_5_796 VPWR VGND sg13g2_decap_8
XFILLER_45_1013 VPWR VGND sg13g2_decap_8
XFILLER_4_295 VPWR VGND sg13g2_decap_8
XFILLER_1_980 VPWR VGND sg13g2_decap_8
X_3120_ _2434_ net987 _0357_ VPWR VGND sg13g2_nor2_1
XFILLER_0_490 VPWR VGND sg13g2_decap_8
X_3051_ ppwm_i.u_ppwm.u_mem.memory\[88\] net792 net794 _2405_ VPWR VGND sg13g2_nor3_1
XFILLER_36_612 VPWR VGND sg13g2_decap_4
XFILLER_36_667 VPWR VGND sg13g2_decap_4
XFILLER_23_317 VPWR VGND sg13g2_decap_8
XFILLER_16_380 VPWR VGND sg13g2_fill_1
X_3953_ net841 VPWR _1005_ VGND ppwm_i.u_ppwm.u_mem.memory\[97\] net648 sg13g2_o21ai_1
X_2904_ _2258_ net1031 VPWR VGND sg13g2_inv_2
X_3884_ VGND VPWR _2192_ net649 _0161_ _0970_ sg13g2_a21oi_1
X_2835_ VPWR _2189_ net903 VGND sg13g2_inv_1
X_5554_ net219 VGND VPWR net1149 falu_i.falutop.alu_data_in\[0\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_4505_ VPWR VGND _1426_ _1455_ _1425_ net616 _1456_ _1413_ sg13g2_a221oi_1
X_5485_ net315 VGND VPWR net998 falu_i.falutop.i2c_inst.sda_o clknet_leaf_6_clk sg13g2_dfrbpq_1
X_4436_ VGND VPWR _1233_ _1327_ _1388_ net640 sg13g2_a21oi_1
X_4367_ _1219_ VPWR _1320_ VGND net615 _1319_ sg13g2_o21ai_1
X_3318_ _0498_ net788 net613 VPWR VGND sg13g2_xnor2_1
Xfanout569 _0814_ net569 VPWR VGND sg13g2_buf_8
X_4298_ _1234_ _1250_ _1251_ VPWR VGND sg13g2_and2_1
XFILLER_39_461 VPWR VGND sg13g2_decap_4
X_3249_ _0442_ net1120 _0440_ VPWR VGND sg13g2_xnor2_1
XFILLER_41_114 VPWR VGND sg13g2_decap_4
XFILLER_41_103 VPWR VGND sg13g2_decap_8
X_5453__74 VPWR VGND net74 sg13g2_tiehi
XFILLER_25_78 VPWR VGND sg13g2_fill_2
XFILLER_10_501 VPWR VGND sg13g2_fill_1
XFILLER_23_884 VPWR VGND sg13g2_decap_8
XFILLER_29_1019 VPWR VGND sg13g2_decap_8
XFILLER_49_269 VPWR VGND sg13g2_decap_8
XFILLER_49_258 VPWR VGND sg13g2_decap_8
XFILLER_46_965 VPWR VGND sg13g2_decap_8
XFILLER_45_442 VPWR VGND sg13g2_decap_8
XFILLER_18_678 VPWR VGND sg13g2_decap_4
XFILLER_32_114 VPWR VGND sg13g2_decap_8
XFILLER_33_626 VPWR VGND sg13g2_fill_2
X_5514__229 VPWR VGND net229 sg13g2_tiehi
XFILLER_14_873 VPWR VGND sg13g2_decap_8
X_5484__317 VPWR VGND net317 sg13g2_tiehi
X_5270_ net156 VGND VPWR net925 ppwm_i.u_ppwm.u_pwm.cmp_value\[8\] clknet_leaf_15_clk
+ sg13g2_dfrbpq_1
X_4221_ net780 _2151_ _1188_ VPWR VGND sg13g2_nor2_1
X_4152_ net1005 net413 _1103_ _0256_ VPWR VGND sg13g2_mux2_1
XFILLER_49_770 VPWR VGND sg13g2_decap_8
X_4083_ _1087_ _1085_ _1086_ VPWR VGND sg13g2_nand2_1
X_3103_ net1014 _0344_ _0345_ VPWR VGND sg13g2_nor2_1
XFILLER_37_943 VPWR VGND sg13g2_decap_8
X_3034_ VPWR VGND _2387_ net786 _2385_ _2383_ _2388_ _2384_ sg13g2_a221oi_1
XFILLER_36_464 VPWR VGND sg13g2_decap_4
X_4985_ net774 VPWR _1928_ VGND falu_i.falutop.div_inst.rem\[1\] falu_i.falutop.div_inst.rem\[0\]
+ sg13g2_o21ai_1
X_3936_ VGND VPWR _2173_ net646 _0187_ _0996_ sg13g2_a21oi_1
XFILLER_20_832 VPWR VGND sg13g2_decap_8
XFILLER_32_670 VPWR VGND sg13g2_fill_2
X_3867_ net825 VPWR _0962_ VGND net443 net657 sg13g2_o21ai_1
XFILLER_31_180 VPWR VGND sg13g2_fill_2
X_3798_ VGND VPWR _2221_ net653 _0118_ _0927_ sg13g2_a21oi_1
X_2818_ VPWR _2172_ net502 VGND sg13g2_inv_1
X_5537_ net84 VGND VPWR net1058 falu_i.falutop.i2c_inst.result\[1\] clknet_leaf_39_clk
+ sg13g2_dfrbpq_1
X_5468_ net349 VGND VPWR _0227_ falu_i.falutop.div_inst.start clknet_leaf_43_clk sg13g2_dfrbpq_2
X_5399_ net254 VGND VPWR _0158_ ppwm_i.u_ppwm.u_mem.memory\[58\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_4419_ _1371_ _1332_ _1286_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_910 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_4
XFILLER_28_987 VPWR VGND sg13g2_decap_8
XFILLER_43_968 VPWR VGND sg13g2_decap_8
XFILLER_14_136 VPWR VGND sg13g2_decap_8
XFILLER_35_1012 VPWR VGND sg13g2_decap_8
XFILLER_11_810 VPWR VGND sg13g2_fill_2
XFILLER_11_832 VPWR VGND sg13g2_decap_8
XFILLER_23_692 VPWR VGND sg13g2_fill_1
XFILLER_22_180 VPWR VGND sg13g2_fill_1
XFILLER_28_8 VPWR VGND sg13g2_fill_2
XFILLER_19_954 VPWR VGND sg13g2_decap_8
XFILLER_45_250 VPWR VGND sg13g2_fill_1
XFILLER_18_464 VPWR VGND sg13g2_decap_4
XFILLER_18_486 VPWR VGND sg13g2_decap_8
XFILLER_45_294 VPWR VGND sg13g2_fill_1
XFILLER_33_434 VPWR VGND sg13g2_fill_2
X_4770_ _1717_ net1037 _1716_ VPWR VGND sg13g2_xnor2_1
XFILLER_14_692 VPWR VGND sg13g2_decap_4
XFILLER_20_128 VPWR VGND sg13g2_fill_1
X_3721_ VGND VPWR net581 _0776_ _0880_ _0879_ sg13g2_a21oi_1
XFILLER_9_184 VPWR VGND sg13g2_fill_2
X_3652_ net608 ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] _0818_ VPWR VGND sg13g2_xor2_1
X_3583_ _0633_ _0694_ _0753_ VPWR VGND sg13g2_nor2_1
X_5322_ net57 VGND VPWR _0081_ ppwm_i.u_ppwm.pwm_value\[9\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_47_0 VPWR VGND sg13g2_decap_8
X_5253_ net189 VGND VPWR _0015_ falu_i.falutop.i2c_inst.data_in\[11\] clknet_leaf_6_clk
+ sg13g2_dfrbpq_1
X_4204_ _1174_ VPWR _1175_ VGND net549 net567 sg13g2_o21ai_1
X_5184_ net1101 net730 net618 _0324_ VPWR VGND sg13g2_mux2_1
X_4135_ net797 _1135_ _0247_ VPWR VGND sg13g2_nor2_1
XFILLER_3_92 VPWR VGND sg13g2_decap_8
XFILLER_28_217 VPWR VGND sg13g2_decap_8
XFILLER_28_228 VPWR VGND sg13g2_decap_4
X_4066_ net871 net777 net684 _0235_ VPWR VGND sg13g2_mux2_1
X_3017_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[48\] net692 _2371_ net708 sg13g2_a21oi_1
X_5495__287 VPWR VGND net287 sg13g2_tiehi
XFILLER_25_946 VPWR VGND sg13g2_decap_8
X_4968_ _1911_ _1909_ _1910_ VPWR VGND sg13g2_xnor2_1
XFILLER_11_128 VPWR VGND sg13g2_fill_1
XFILLER_12_629 VPWR VGND sg13g2_decap_4
X_3919_ net834 VPWR _0988_ VGND net886 net647 sg13g2_o21ai_1
X_4899_ _1820_ VPWR _1843_ VGND _1799_ _1821_ sg13g2_o21ai_1
XFILLER_20_651 VPWR VGND sg13g2_decap_8
XFILLER_16_902 VPWR VGND sg13g2_decap_8
XFILLER_43_721 VPWR VGND sg13g2_decap_4
XFILLER_43_776 VPWR VGND sg13g2_fill_2
XFILLER_42_242 VPWR VGND sg13g2_decap_8
XFILLER_16_979 VPWR VGND sg13g2_decap_8
XFILLER_30_415 VPWR VGND sg13g2_fill_2
XFILLER_11_651 VPWR VGND sg13g2_fill_1
X_5253__189 VPWR VGND net189 sg13g2_tiehi
XFILLER_7_655 VPWR VGND sg13g2_decap_4
XFILLER_6_121 VPWR VGND sg13g2_decap_8
XFILLER_40_7 VPWR VGND sg13g2_fill_2
XFILLER_3_861 VPWR VGND sg13g2_decap_8
Xheichips25_tiny_wrapper_19 VPWR VGND uio_out[3] sg13g2_tielo
XFILLER_19_4 VPWR VGND sg13g2_decap_4
XFILLER_19_751 VPWR VGND sg13g2_decap_8
XFILLER_19_773 VPWR VGND sg13g2_fill_2
X_4822_ _1768_ _1765_ _1767_ VPWR VGND sg13g2_nand2_1
X_4753_ _1698_ _1697_ _1692_ _1700_ VPWR VGND sg13g2_a21o_1
X_3704_ _0864_ _2237_ net601 VPWR VGND sg13g2_xnor2_1
XFILLER_30_993 VPWR VGND sg13g2_decap_8
X_4684_ _1631_ _1392_ _1632_ VPWR VGND sg13g2_xor2_1
X_3635_ net585 _0719_ _0802_ VPWR VGND sg13g2_nor2_1
X_3566_ net609 _0719_ _0737_ VPWR VGND sg13g2_nor2_1
X_5305_ net223 VGND VPWR net387 ppwm_i.u_ppwm.u_ex.state_q\[1\] clknet_leaf_20_clk
+ sg13g2_dfrbpq_1
X_3497_ net575 _0670_ _0671_ VPWR VGND sg13g2_and2_1
X_5236_ VGND VPWR net626 _2142_ _0341_ _2141_ sg13g2_a21oi_1
X_5167_ net1148 net620 _2102_ VPWR VGND sg13g2_nor2_1
X_5098_ VGND VPWR _1985_ _2002_ _2038_ _2001_ sg13g2_a21oi_1
X_4118_ _1120_ falu_i.falutop.div_inst.b1\[2\] falu_i.falutop.div_inst.acc\[2\] VPWR
+ VGND sg13g2_xnor2_1
X_4049_ VGND VPWR _2441_ _0901_ _1071_ _1057_ sg13g2_a21oi_1
XFILLER_37_581 VPWR VGND sg13g2_decap_8
XFILLER_25_721 VPWR VGND sg13g2_decap_8
XFILLER_24_242 VPWR VGND sg13g2_fill_1
XFILLER_9_909 VPWR VGND sg13g2_decap_8
XFILLER_12_415 VPWR VGND sg13g2_decap_8
XFILLER_12_426 VPWR VGND sg13g2_fill_1
XFILLER_3_113 VPWR VGND sg13g2_fill_2
XFILLER_3_157 VPWR VGND sg13g2_fill_2
XFILLER_0_820 VPWR VGND sg13g2_decap_8
Xhold8 falu_i.falutop.div_inst.done VPWR VGND net380 sg13g2_dlygate4sd3_1
XFILLER_0_897 VPWR VGND sg13g2_decap_8
XFILLER_48_879 VPWR VGND sg13g2_decap_8
XFILLER_15_220 VPWR VGND sg13g2_fill_2
XFILLER_43_540 VPWR VGND sg13g2_decap_8
XFILLER_31_735 VPWR VGND sg13g2_fill_2
XFILLER_30_256 VPWR VGND sg13g2_fill_2
XFILLER_12_993 VPWR VGND sg13g2_decap_8
Xhold408 ppwm_i.u_ppwm.u_pwm.counter\[5\] VPWR VGND net1060 sg13g2_dlygate4sd3_1
XFILLER_8_986 VPWR VGND sg13g2_decap_8
XFILLER_7_474 VPWR VGND sg13g2_decap_8
X_3420_ VPWR VGND ppwm_i.u_ppwm.pwm_value\[7\] _0597_ _2260_ ppwm_i.u_ppwm.pwm_value\[8\]
+ _0598_ _2259_ sg13g2_a221oi_1
Xhold419 falu_i.falutop.i2c_inst.result\[14\] VPWR VGND net1071 sg13g2_dlygate4sd3_1
X_3351_ _0517_ VPWR _0529_ VGND _0518_ _0528_ sg13g2_o21ai_1
X_5561__141 VPWR VGND net141 sg13g2_tiehi
X_5346__360 VPWR VGND net360 sg13g2_tiehi
X_3282_ VPWR VGND ppwm_i.u_ppwm.u_pwm.counter\[3\] _0464_ _2285_ ppwm_i.u_ppwm.u_pwm.counter\[4\]
+ _0465_ _2284_ sg13g2_a221oi_1
X_5021_ _1933_ _1962_ _1963_ VPWR VGND sg13g2_nor2_1
XFILLER_24_2 VPWR VGND sg13g2_fill_1
XFILLER_38_345 VPWR VGND sg13g2_decap_4
XFILLER_0_1002 VPWR VGND sg13g2_decap_8
XFILLER_47_890 VPWR VGND sg13g2_decap_8
X_4805_ net713 net766 _1751_ VPWR VGND sg13g2_and2_1
XFILLER_10_908 VPWR VGND sg13g2_decap_8
XFILLER_22_768 VPWR VGND sg13g2_decap_8
X_2997_ _2351_ net690 ppwm_i.u_ppwm.u_mem.memory\[93\] net702 ppwm_i.u_ppwm.u_mem.memory\[107\]
+ VPWR VGND sg13g2_a22oi_1
X_4736_ _1683_ net746 net748 VPWR VGND sg13g2_nand2_1
XFILLER_30_790 VPWR VGND sg13g2_decap_4
X_4667_ _1615_ _1327_ _1215_ _1324_ _1216_ VPWR VGND sg13g2_a22oi_1
X_3618_ net576 _0784_ _0786_ VPWR VGND _0785_ sg13g2_nand3b_1
X_4598_ net754 net726 net566 _1547_ VPWR VGND sg13g2_mux2_1
X_3549_ _0721_ _0720_ _0622_ _0678_ net571 VPWR VGND sg13g2_a22oi_1
X_5219_ _2129_ falu_i.falutop.data_in\[9\] _2130_ VPWR VGND sg13g2_xor2_1
XFILLER_44_348 VPWR VGND sg13g2_decap_8
XFILLER_13_702 VPWR VGND sg13g2_fill_1
XFILLER_12_256 VPWR VGND sg13g2_fill_2
XFILLER_5_923 VPWR VGND sg13g2_decap_8
XFILLER_4_433 VPWR VGND sg13g2_fill_2
XFILLER_4_466 VPWR VGND sg13g2_fill_1
XFILLER_4_488 VPWR VGND sg13g2_fill_2
XFILLER_47_120 VPWR VGND sg13g2_fill_2
X_5556__210 VPWR VGND net210 sg13g2_tiehi
XFILLER_36_827 VPWR VGND sg13g2_decap_4
XFILLER_47_186 VPWR VGND sg13g2_fill_2
XFILLER_35_337 VPWR VGND sg13g2_decap_8
X_2920_ VPWR _2274_ net1094 VGND sg13g2_inv_1
XFILLER_16_595 VPWR VGND sg13g2_decap_8
X_2851_ VPWR _2205_ net854 VGND sg13g2_inv_1
XFILLER_12_790 VPWR VGND sg13g2_fill_2
X_5570_ net64 VGND VPWR net1082 falu_i.falutop.div_inst.b\[0\] clknet_leaf_4_clk sg13g2_dfrbpq_1
XFILLER_31_598 VPWR VGND sg13g2_fill_2
X_4521_ _1469_ _1466_ _1471_ VPWR VGND sg13g2_xor2_1
Xhold205 _0290_ VPWR VGND net857 sg13g2_dlygate4sd3_1
X_4452_ net776 falu_i.falutop.data_in\[7\] _1404_ VPWR VGND sg13g2_xor2_1
Xhold216 ppwm_i.u_ppwm.u_mem.memory\[0\] VPWR VGND net868 sg13g2_dlygate4sd3_1
X_3403_ _0581_ ppwm_i.u_ppwm.u_ex.reg_value_q\[9\] _2258_ VPWR VGND sg13g2_nand2_1
Xhold238 _0166_ VPWR VGND net890 sg13g2_dlygate4sd3_1
Xhold227 falu_i.falutop.div_inst.acc\[8\] VPWR VGND net879 sg13g2_dlygate4sd3_1
Xhold249 falu_i.falutop.i2c_inst.data_in\[1\] VPWR VGND net901 sg13g2_dlygate4sd3_1
X_4383_ _1335_ _1333_ _1331_ _1336_ VPWR VGND sg13g2_a21o_1
X_3334_ _0512_ VPWR _0513_ VGND _2253_ _0510_ sg13g2_o21ai_1
Xfanout718 net719 net718 VPWR VGND sg13g2_buf_8
Xfanout729 falu_i.falutop.alu_data_in\[12\] net729 VPWR VGND sg13g2_buf_8
Xfanout707 _2295_ net707 VPWR VGND sg13g2_buf_8
X_3265_ net796 _0451_ _0452_ _0060_ VPWR VGND sg13g2_nor3_1
X_5311__79 VPWR VGND net79 sg13g2_tiehi
X_5004_ _1945_ VPWR _1946_ VGND _1906_ _1911_ sg13g2_o21ai_1
XFILLER_39_687 VPWR VGND sg13g2_fill_1
XFILLER_27_827 VPWR VGND sg13g2_fill_2
X_3196_ net1049 _0402_ net863 _0407_ VPWR VGND sg13g2_nand3_1
X_5500__275 VPWR VGND net275 sg13g2_tiehi
XFILLER_14_14 VPWR VGND sg13g2_decap_4
X_4719_ VGND VPWR _2297_ net565 _1666_ _1665_ sg13g2_a21oi_1
XFILLER_5_219 VPWR VGND sg13g2_decap_8
XFILLER_2_904 VPWR VGND sg13g2_decap_8
XFILLER_30_79 VPWR VGND sg13g2_fill_1
XFILLER_1_436 VPWR VGND sg13g2_decap_8
XFILLER_1_447 VPWR VGND sg13g2_decap_4
XFILLER_18_816 VPWR VGND sg13g2_decap_8
XFILLER_29_164 VPWR VGND sg13g2_fill_1
XFILLER_26_860 VPWR VGND sg13g2_decap_8
XFILLER_41_874 VPWR VGND sg13g2_fill_1
XFILLER_13_554 VPWR VGND sg13g2_fill_2
XFILLER_9_536 VPWR VGND sg13g2_decap_4
XFILLER_5_731 VPWR VGND sg13g2_fill_1
X_3050_ VGND VPWR _2403_ _2404_ _2397_ _2394_ sg13g2_a21oi_2
XFILLER_49_985 VPWR VGND sg13g2_decap_8
X_3952_ VGND VPWR _2167_ net677 _0195_ _1004_ sg13g2_a21oi_1
X_2903_ VPWR _2257_ net793 VGND sg13g2_inv_1
X_3883_ net839 VPWR _0970_ VGND net474 net649 sg13g2_o21ai_1
XFILLER_32_885 VPWR VGND sg13g2_fill_1
X_2834_ VPWR _2188_ net889 VGND sg13g2_inv_1
XFILLER_31_384 VPWR VGND sg13g2_decap_4
X_5553_ net227 VGND VPWR _0312_ falu_i.falutop.div_inst.b\[7\] clknet_leaf_3_clk sg13g2_dfrbpq_1
X_4504_ _1450_ VPWR _1455_ VGND _1451_ _1454_ sg13g2_o21ai_1
X_5484_ net317 VGND VPWR net909 falu_i.falutop.data_in\[15\] clknet_leaf_6_clk sg13g2_dfrbpq_1
X_4435_ _1387_ _1385_ net631 _1375_ _1373_ VPWR VGND sg13g2_a22oi_1
X_4366_ net772 net771 _1279_ _1319_ VPWR VGND sg13g2_nor3_2
X_3317_ _0497_ net788 net613 VPWR VGND sg13g2_nand2_1
X_4297_ _1248_ _1239_ _1250_ VPWR VGND sg13g2_xor2_1
X_3248_ _0440_ net1140 _0054_ VPWR VGND sg13g2_nor2_1
XFILLER_27_602 VPWR VGND sg13g2_fill_2
X_3179_ net810 VPWR _0395_ VGND ppwm_i.u_ppwm.pwm_value\[8\] net682 sg13g2_o21ai_1
XFILLER_39_495 VPWR VGND sg13g2_decap_8
XFILLER_26_112 VPWR VGND sg13g2_fill_1
XFILLER_23_863 VPWR VGND sg13g2_decap_8
XFILLER_22_395 VPWR VGND sg13g2_fill_2
XFILLER_49_237 VPWR VGND sg13g2_decap_8
X_5403__246 VPWR VGND net246 sg13g2_tiehi
XFILLER_46_944 VPWR VGND sg13g2_decap_8
XFILLER_33_638 VPWR VGND sg13g2_decap_4
XFILLER_14_852 VPWR VGND sg13g2_decap_8
XFILLER_41_682 VPWR VGND sg13g2_decap_8
X_4220_ VGND VPWR net606 _1186_ _0280_ _1187_ sg13g2_a21oi_1
X_4151_ VPWR _0255_ net480 VGND sg13g2_inv_1
X_4082_ _1086_ _0343_ falu_i.falutop.i2c_inst.result\[2\] _2445_ falu_i.falutop.i2c_inst.result\[1\]
+ VPWR VGND sg13g2_a22oi_1
X_3102_ _0344_ _2433_ net1046 VPWR VGND sg13g2_nand2_2
X_3033_ VPWR VGND _2226_ _2386_ net688 _2216_ _2387_ net700 sg13g2_a221oi_1
XFILLER_36_421 VPWR VGND sg13g2_decap_4
XFILLER_36_443 VPWR VGND sg13g2_decap_8
XFILLER_37_999 VPWR VGND sg13g2_decap_8
X_4984_ VGND VPWR _1927_ _1926_ _1923_ sg13g2_or2_1
XFILLER_24_638 VPWR VGND sg13g2_decap_8
X_3935_ net836 VPWR _0996_ VGND ppwm_i.u_ppwm.u_mem.memory\[88\] net646 sg13g2_o21ai_1
XFILLER_20_811 VPWR VGND sg13g2_decap_8
X_3866_ VGND VPWR _2198_ net657 _0152_ _0961_ sg13g2_a21oi_1
XFILLER_20_888 VPWR VGND sg13g2_decap_8
X_3797_ net827 VPWR _0927_ VGND net898 net653 sg13g2_o21ai_1
X_2817_ VPWR _2171_ net957 VGND sg13g2_inv_1
X_5536_ net96 VGND VPWR net1023 falu_i.falutop.i2c_inst.result\[0\] clknet_leaf_38_clk
+ sg13g2_dfrbpq_1
X_5467_ net353 VGND VPWR _0226_ falu_i.falutop.i2c_inst.counter\[4\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_4418_ _1365_ VPWR _1370_ VGND _1289_ _1369_ sg13g2_o21ai_1
X_5398_ net256 VGND VPWR net558 ppwm_i.u_ppwm.u_mem.memory\[57\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_4349_ falu_i.falutop.alu_inst.op\[1\] falu_i.falutop.alu_inst.op\[0\] _1302_ VPWR
+ VGND sg13g2_nor2_1
XFILLER_28_966 VPWR VGND sg13g2_decap_8
XFILLER_27_487 VPWR VGND sg13g2_decap_8
XFILLER_43_947 VPWR VGND sg13g2_decap_8
XFILLER_42_457 VPWR VGND sg13g2_fill_1
XFILLER_11_888 VPWR VGND sg13g2_decap_8
XFILLER_10_398 VPWR VGND sg13g2_fill_2
X_5286__125 VPWR VGND net125 sg13g2_tiehi
XFILLER_19_933 VPWR VGND sg13g2_decap_8
XFILLER_46_763 VPWR VGND sg13g2_fill_2
X_5438__139 VPWR VGND net139 sg13g2_tiehi
XFILLER_34_969 VPWR VGND sg13g2_decap_8
X_3720_ net578 VPWR _0879_ VGND ppwm_i.u_ppwm.pwm_value\[7\] net583 sg13g2_o21ai_1
XFILLER_42_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_40_clk clknet_3_1__leaf_clk clknet_leaf_40_clk VPWR VGND sg13g2_buf_8
X_3651_ VGND VPWR net582 _0640_ _0817_ _0816_ sg13g2_a21oi_1
X_3582_ _0751_ VPWR _0752_ VGND _0746_ _0749_ sg13g2_o21ai_1
X_5321_ net59 VGND VPWR _0080_ ppwm_i.u_ppwm.pwm_value\[8\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_6_892 VPWR VGND sg13g2_decap_8
XFILLER_5_391 VPWR VGND sg13g2_decap_4
X_5252_ net191 VGND VPWR _0014_ falu_i.falutop.i2c_inst.data_in\[10\] clknet_leaf_7_clk
+ sg13g2_dfrbpq_1
X_4203_ _1174_ net567 _1173_ VPWR VGND sg13g2_nand2_1
X_5183_ net1122 net735 net618 _0323_ VPWR VGND sg13g2_mux2_1
X_4134_ VGND VPWR net779 _1102_ _1135_ net633 sg13g2_a21oi_1
XFILLER_37_741 VPWR VGND sg13g2_decap_8
XFILLER_3_1022 VPWR VGND sg13g2_decap_8
X_4065_ net850 falu_i.falutop.data_in\[6\] net684 _0234_ VPWR VGND sg13g2_mux2_1
X_3016_ ppwm_i.u_ppwm.u_mem.memory\[41\] net688 _2370_ VPWR VGND sg13g2_and2_1
XFILLER_25_925 VPWR VGND sg13g2_decap_8
X_5356__340 VPWR VGND net340 sg13g2_tiehi
XFILLER_24_468 VPWR VGND sg13g2_fill_1
XFILLER_40_939 VPWR VGND sg13g2_decap_8
X_4967_ _1910_ _1859_ _2304_ _1858_ _1751_ VPWR VGND sg13g2_a22oi_1
X_3918_ VGND VPWR _2179_ net669 _0178_ _0987_ sg13g2_a21oi_1
X_4898_ VGND VPWR _1792_ _1796_ _1842_ _1798_ sg13g2_a21oi_1
XFILLER_22_25 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_31_clk clknet_3_7__leaf_clk clknet_leaf_31_clk VPWR VGND sg13g2_buf_8
X_3849_ net831 VPWR _0953_ VGND net860 net664 sg13g2_o21ai_1
X_5519_ net206 VGND VPWR _0278_ falu_i.falutop.div_inst.rem\[6\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_229 VPWR VGND sg13g2_fill_2
XFILLER_28_730 VPWR VGND sg13g2_decap_4
XFILLER_42_221 VPWR VGND sg13g2_fill_1
XFILLER_15_413 VPWR VGND sg13g2_decap_4
XFILLER_16_958 VPWR VGND sg13g2_decap_8
XFILLER_15_457 VPWR VGND sg13g2_decap_8
XFILLER_15_468 VPWR VGND sg13g2_fill_1
XFILLER_43_799 VPWR VGND sg13g2_decap_8
XFILLER_15_479 VPWR VGND sg13g2_decap_4
XFILLER_24_991 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_22_clk clknet_3_4__leaf_clk clknet_leaf_22_clk VPWR VGND sg13g2_buf_8
XFILLER_30_449 VPWR VGND sg13g2_fill_2
XFILLER_7_634 VPWR VGND sg13g2_decap_4
XFILLER_7_601 VPWR VGND sg13g2_fill_2
XFILLER_11_685 VPWR VGND sg13g2_decap_8
XFILLER_6_133 VPWR VGND sg13g2_decap_4
XFILLER_3_840 VPWR VGND sg13g2_decap_8
XFILLER_46_560 VPWR VGND sg13g2_fill_1
XFILLER_34_722 VPWR VGND sg13g2_fill_1
X_4821_ _1764_ _1763_ _1758_ _1767_ VPWR VGND sg13g2_a21o_1
XFILLER_33_243 VPWR VGND sg13g2_decap_8
XFILLER_15_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk clknet_leaf_13_clk VPWR VGND sg13g2_buf_8
X_4752_ _1697_ _1698_ _1692_ _1699_ VPWR VGND sg13g2_nand3_1
X_3703_ VPWR VGND _0863_ net795 _0860_ _2238_ _0087_ net569 sg13g2_a221oi_1
X_4683_ VGND VPWR _1224_ _1227_ _1631_ _1630_ sg13g2_a21oi_1
XFILLER_30_972 VPWR VGND sg13g2_decap_8
X_3634_ VGND VPWR _0798_ _0799_ _0801_ _0800_ sg13g2_a21oi_1
X_3565_ net574 _0733_ _0734_ _0735_ _0736_ VPWR VGND sg13g2_nor4_1
X_5304_ net95 VGND VPWR net982 ppwm_i.u_ppwm.u_ex.state_q\[0\] clknet_leaf_19_clk
+ sg13g2_dfrbpq_1
X_3496_ _0670_ _0668_ _0669_ VPWR VGND sg13g2_nand2_1
X_5235_ _2142_ falu_i.falutop.data_in\[13\] _2140_ VPWR VGND sg13g2_xnor2_1
XFILLER_25_1023 VPWR VGND sg13g2_decap_4
X_5166_ VPWR _0312_ net1075 VGND sg13g2_inv_1
XFILLER_29_516 VPWR VGND sg13g2_fill_1
XFILLER_29_505 VPWR VGND sg13g2_decap_8
X_5097_ _2037_ _2019_ _2036_ VPWR VGND sg13g2_xnor2_1
X_4117_ _1116_ VPWR _1119_ VGND _1117_ _1118_ sg13g2_o21ai_1
XFILLER_17_47 VPWR VGND sg13g2_fill_1
X_4048_ net797 _1070_ _0225_ VPWR VGND sg13g2_nor2_1
XFILLER_24_254 VPWR VGND sg13g2_fill_1
XFILLER_21_994 VPWR VGND sg13g2_decap_8
XFILLER_4_648 VPWR VGND sg13g2_fill_1
XFILLER_48_814 VPWR VGND sg13g2_fill_1
XFILLER_0_876 VPWR VGND sg13g2_decap_8
Xhold9 ppwm_i.u_ppwm.u_pwm.cmp_value\[0\] VPWR VGND net381 sg13g2_dlygate4sd3_1
XFILLER_48_858 VPWR VGND sg13g2_decap_8
XFILLER_16_744 VPWR VGND sg13g2_decap_8
XFILLER_31_725 VPWR VGND sg13g2_fill_1
XFILLER_12_972 VPWR VGND sg13g2_decap_8
XFILLER_8_965 VPWR VGND sg13g2_decap_8
Xhold409 _0039_ VPWR VGND net1061 sg13g2_dlygate4sd3_1
XFILLER_7_453 VPWR VGND sg13g2_fill_2
XFILLER_7_486 VPWR VGND sg13g2_decap_8
XFILLER_48_1012 VPWR VGND sg13g2_decap_8
X_3350_ VPWR VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] _0527_ _2245_ net782 _0528_
+ _2244_ sg13g2_a221oi_1
X_5308__85 VPWR VGND net85 sg13g2_tiehi
XFILLER_3_681 VPWR VGND sg13g2_fill_2
X_5323__55 VPWR VGND net55 sg13g2_tiehi
X_5020_ _1962_ _1934_ _1960_ VPWR VGND sg13g2_xnor2_1
X_3281_ VPWR VGND _0462_ _0463_ _0461_ _2278_ _0464_ ppwm_i.u_ppwm.u_pwm.cmp_value\[3\]
+ sg13g2_a221oi_1
XFILLER_39_814 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk clknet_leaf_2_clk VPWR VGND sg13g2_buf_8
XFILLER_39_847 VPWR VGND sg13g2_fill_2
X_4804_ _1750_ net732 net753 VPWR VGND sg13g2_nand2_1
X_2996_ _2348_ _2349_ _2347_ _2350_ VPWR VGND sg13g2_nand3_1
X_4735_ VGND VPWR _1682_ _1625_ _1623_ sg13g2_or2_1
X_4666_ VPWR VGND _1217_ _1363_ _1383_ _1214_ _1614_ _1319_ sg13g2_a221oi_1
X_3617_ _0782_ _0783_ _0785_ VPWR VGND sg13g2_nor2b_1
X_4597_ _1546_ _1480_ _1544_ VPWR VGND sg13g2_xnor2_1
X_3548_ _0700_ _0719_ net609 _0720_ VPWR VGND sg13g2_mux2_1
X_3479_ VGND VPWR net609 _0626_ _0654_ _0653_ sg13g2_a21oi_1
X_5218_ _2129_ net775 falu_i.falutop.data_in\[8\] VPWR VGND sg13g2_nand2_1
X_5149_ _2087_ falu_i.falutop.div_inst.rem\[7\] _2086_ VPWR VGND sg13g2_xnor2_1
XFILLER_28_35 VPWR VGND sg13g2_fill_1
XFILLER_44_327 VPWR VGND sg13g2_fill_1
XFILLER_40_511 VPWR VGND sg13g2_decap_8
XFILLER_13_736 VPWR VGND sg13g2_decap_8
XFILLER_13_758 VPWR VGND sg13g2_decap_8
XFILLER_13_769 VPWR VGND sg13g2_fill_1
XFILLER_21_791 VPWR VGND sg13g2_decap_8
XFILLER_5_902 VPWR VGND sg13g2_decap_8
XFILLER_5_979 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_688 VPWR VGND sg13g2_decap_4
X_5517__217 VPWR VGND net217 sg13g2_tiehi
XFILLER_43_360 VPWR VGND sg13g2_decap_8
X_2850_ VPWR _2204_ net893 VGND sg13g2_inv_1
X_5413__226 VPWR VGND net226 sg13g2_tiehi
XFILLER_15_1022 VPWR VGND sg13g2_decap_8
X_4520_ _1466_ _1469_ _1470_ VPWR VGND sg13g2_nor2_1
X_4451_ net818 VPWR _1403_ VGND net1057 net628 sg13g2_o21ai_1
Xhold206 falu_i.falutop.i2c_inst.data_in\[11\] VPWR VGND net858 sg13g2_dlygate4sd3_1
Xhold217 falu_i.falutop.i2c_inst.data_in\[5\] VPWR VGND net869 sg13g2_dlygate4sd3_1
X_3402_ ppwm_i.u_ppwm.global_counter\[17\] _2236_ _0579_ _0580_ VPWR VGND sg13g2_a21o_1
Xhold228 _1213_ VPWR VGND net880 sg13g2_dlygate4sd3_1
Xhold239 falu_i.falutop.div_inst.b\[2\] VPWR VGND net891 sg13g2_dlygate4sd3_1
X_4382_ net726 _1334_ _1335_ VPWR VGND sg13g2_nor2_1
Xfanout708 _2256_ net708 VPWR VGND sg13g2_buf_8
X_3333_ _0479_ _0511_ _0512_ VPWR VGND sg13g2_nor2_1
Xfanout719 net720 net719 VPWR VGND sg13g2_buf_1
X_3264_ _2262_ _0449_ _0452_ VPWR VGND sg13g2_nor2_2
X_5003_ VPWR _1945_ _1944_ VGND sg13g2_inv_1
X_3195_ _0406_ net863 ppwm_i.u_ppwm.u_pwm.counter\[2\] VPWR VGND sg13g2_nand2_1
XFILLER_38_176 VPWR VGND sg13g2_decap_8
XFILLER_10_717 VPWR VGND sg13g2_fill_1
X_2979_ _2333_ net697 _2175_ net702 _2161_ VPWR VGND sg13g2_a22oi_1
X_4718_ net747 net565 _1665_ VPWR VGND sg13g2_nor2_1
X_4649_ _1597_ _1595_ _1596_ VPWR VGND sg13g2_nand2_1
X_5456__62 VPWR VGND net62 sg13g2_tiehi
XFILLER_44_113 VPWR VGND sg13g2_fill_2
XFILLER_9_504 VPWR VGND sg13g2_decap_4
XFILLER_49_964 VPWR VGND sg13g2_decap_8
XFILLER_48_463 VPWR VGND sg13g2_fill_2
X_5296__105 VPWR VGND net105 sg13g2_tiehi
XFILLER_36_636 VPWR VGND sg13g2_fill_2
XFILLER_24_809 VPWR VGND sg13g2_decap_8
X_3951_ net840 VPWR _1004_ VGND net556 net677 sg13g2_o21ai_1
XFILLER_17_883 VPWR VGND sg13g2_decap_8
XFILLER_44_691 VPWR VGND sg13g2_decap_4
X_2902_ VPWR _2256_ net789 VGND sg13g2_inv_1
XFILLER_16_371 VPWR VGND sg13g2_decap_8
XFILLER_43_190 VPWR VGND sg13g2_fill_2
X_3882_ VGND VPWR _2192_ net676 _0160_ _0969_ sg13g2_a21oi_1
XFILLER_31_330 VPWR VGND sg13g2_fill_2
X_2833_ VPWR _2187_ net904 VGND sg13g2_inv_1
XFILLER_31_363 VPWR VGND sg13g2_fill_2
X_5552_ net235 VGND VPWR _0311_ falu_i.falutop.div_inst.a\[7\] clknet_leaf_43_clk
+ sg13g2_dfrbpq_1
X_4503_ VPWR VGND _1453_ _1289_ _1452_ _1284_ _1454_ _1300_ sg13g2_a221oi_1
X_5483_ net319 VGND VPWR net862 falu_i.falutop.data_in\[14\] clknet_leaf_6_clk sg13g2_dfrbpq_2
X_4434_ _1384_ VPWR _1386_ VGND _1231_ _1314_ sg13g2_o21ai_1
X_4365_ VGND VPWR _1318_ _1279_ _1259_ sg13g2_or2_1
X_3316_ VGND VPWR net791 _2418_ _0496_ _0486_ sg13g2_a21oi_1
X_4296_ _1249_ _1239_ _1248_ VPWR VGND sg13g2_nand2_1
X_3247_ net812 VPWR _0441_ VGND net1139 _0439_ sg13g2_o21ai_1
X_5424__196 VPWR VGND net196 sg13g2_tiehi
X_3178_ VGND VPWR _2281_ net683 _0031_ _0394_ sg13g2_a21oi_1
XFILLER_25_14 VPWR VGND sg13g2_fill_2
XFILLER_23_842 VPWR VGND sg13g2_decap_8
XFILLER_22_363 VPWR VGND sg13g2_decap_4
XFILLER_10_558 VPWR VGND sg13g2_fill_2
X_5431__167 VPWR VGND net167 sg13g2_tiehi
X_5366__320 VPWR VGND net320 sg13g2_tiehi
XFILLER_1_201 VPWR VGND sg13g2_fill_1
XFILLER_9_4 VPWR VGND sg13g2_fill_2
XFILLER_49_205 VPWR VGND sg13g2_decap_4
XFILLER_2_18 VPWR VGND sg13g2_fill_2
XFILLER_46_923 VPWR VGND sg13g2_decap_8
XFILLER_45_466 VPWR VGND sg13g2_decap_8
XFILLER_33_628 VPWR VGND sg13g2_fill_1
XFILLER_14_831 VPWR VGND sg13g2_decap_8
XFILLER_32_127 VPWR VGND sg13g2_fill_1
XFILLER_9_301 VPWR VGND sg13g2_fill_2
XFILLER_9_312 VPWR VGND sg13g2_fill_1
XFILLER_13_385 VPWR VGND sg13g2_fill_1
XFILLER_12_1014 VPWR VGND sg13g2_decap_8
X_4150_ _1143_ _1104_ net479 falu_i.falutop.div_inst.b\[0\] net778 VPWR VGND sg13g2_a22oi_1
X_3101_ net1132 falu_i.falutop.i2c_inst.counter\[1\] _0343_ VPWR VGND sg13g2_nor2b_2
X_4081_ _1085_ _2438_ falu_i.falutop.i2c_inst.result\[0\] _2432_ falu_i.falutop.i2c_inst.result\[3\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_49_794 VPWR VGND sg13g2_decap_8
X_3032_ ppwm_i.u_ppwm.u_mem.memory\[5\] net791 net793 _2386_ VPWR VGND sg13g2_nor3_1
XFILLER_48_293 VPWR VGND sg13g2_fill_2
XFILLER_37_978 VPWR VGND sg13g2_decap_8
X_4983_ _1834_ VPWR _1926_ VGND _1924_ _1925_ sg13g2_o21ai_1
XFILLER_23_105 VPWR VGND sg13g2_fill_1
X_3934_ VGND VPWR _2173_ net675 _0186_ _0995_ sg13g2_a21oi_1
X_3865_ net829 VPWR _0961_ VGND ppwm_i.u_ppwm.u_mem.memory\[52\] net665 sg13g2_o21ai_1
XFILLER_20_867 VPWR VGND sg13g2_decap_8
X_2816_ _2170_ net390 VPWR VGND sg13g2_inv_2
X_3796_ VGND VPWR _2222_ net659 _0117_ _0926_ sg13g2_a21oi_1
X_5535_ net104 VGND VPWR _0294_ falu_i.falutop.div_inst.acc\[8\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_5466_ net357 VGND VPWR _0225_ falu_i.falutop.i2c_inst.counter\[3\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_4417_ _1366_ _1368_ _1284_ _1369_ VPWR VGND sg13g2_mux2_1
X_5397_ net258 VGND VPWR net395 ppwm_i.u_ppwm.u_mem.memory\[56\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
X_4348_ _1300_ _1297_ _1288_ _1301_ VPWR VGND sg13g2_mux2_1
X_4279_ net707 _2304_ _1232_ VPWR VGND sg13g2_nor2_2
XFILLER_28_945 VPWR VGND sg13g2_decap_8
XFILLER_43_926 VPWR VGND sg13g2_decap_8
XFILLER_10_333 VPWR VGND sg13g2_fill_2
XFILLER_11_867 VPWR VGND sg13g2_decap_8
XFILLER_22_171 VPWR VGND sg13g2_decap_8
XFILLER_2_521 VPWR VGND sg13g2_decap_8
XFILLER_19_912 VPWR VGND sg13g2_decap_8
XFILLER_19_989 VPWR VGND sg13g2_decap_8
X_5490__301 VPWR VGND net301 sg13g2_tiehi
XFILLER_45_285 VPWR VGND sg13g2_decap_8
XFILLER_34_948 VPWR VGND sg13g2_decap_8
XFILLER_41_491 VPWR VGND sg13g2_decap_8
X_3650_ ppwm_i.u_ppwm.pwm_value\[0\] net582 _0816_ VPWR VGND sg13g2_nor2_1
X_3581_ _0618_ _0750_ _0751_ VPWR VGND sg13g2_nor2_1
XFILLER_9_186 VPWR VGND sg13g2_fill_1
X_5320_ net61 VGND VPWR net1191 ppwm_i.u_ppwm.pwm_value\[7\] clknet_leaf_17_clk sg13g2_dfrbpq_2
XFILLER_6_871 VPWR VGND sg13g2_decap_8
X_5251_ net193 VGND VPWR _0013_ falu_i.falutop.i2c_inst.data_in\[9\] clknet_leaf_37_clk
+ sg13g2_dfrbpq_1
X_4202_ _1173_ _1125_ _1126_ VPWR VGND sg13g2_xnor2_1
X_5182_ VGND VPWR net707 net618 _0322_ _2107_ sg13g2_a21oi_1
X_4133_ _1095_ _1096_ _1134_ VPWR VGND sg13g2_nor2_2
XFILLER_3_1001 VPWR VGND sg13g2_decap_8
X_4064_ net869 falu_i.falutop.data_in\[5\] net684 _0233_ VPWR VGND sg13g2_mux2_1
X_3015_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[20\] net788 net692 ppwm_i.u_ppwm.u_mem.memory\[6\]
+ _2369_ net696 sg13g2_a221oi_1
XFILLER_37_775 VPWR VGND sg13g2_fill_1
XFILLER_25_904 VPWR VGND sg13g2_decap_8
XFILLER_36_296 VPWR VGND sg13g2_decap_8
X_5532__128 VPWR VGND net128 sg13g2_tiehi
X_4966_ _1909_ _1908_ _1907_ VPWR VGND sg13g2_nand2b_1
XFILLER_33_981 VPWR VGND sg13g2_decap_8
X_3917_ net834 VPWR _0987_ VGND ppwm_i.u_ppwm.u_mem.memory\[78\] net669 sg13g2_o21ai_1
X_4897_ _1824_ VPWR _1841_ VGND _1747_ _1825_ sg13g2_o21ai_1
XFILLER_32_491 VPWR VGND sg13g2_decap_8
X_3848_ VGND VPWR _2205_ net643 _0143_ _0952_ sg13g2_a21oi_1
XFILLER_20_675 VPWR VGND sg13g2_decap_8
XFILLER_20_686 VPWR VGND sg13g2_fill_1
X_3779_ net830 VPWR _0918_ VGND ppwm_i.u_ppwm.u_mem.memory\[9\] net662 sg13g2_o21ai_1
X_5518_ net213 VGND VPWR _0277_ falu_i.falutop.div_inst.rem\[5\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_5449_ net91 VGND VPWR net462 ppwm_i.u_ppwm.u_mem.memory\[108\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
XFILLER_16_937 VPWR VGND sg13g2_decap_8
XFILLER_24_970 VPWR VGND sg13g2_decap_8
XFILLER_42_299 VPWR VGND sg13g2_decap_8
XFILLER_7_613 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_decap_4
XFILLER_11_664 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_3_896 VPWR VGND sg13g2_decap_8
XFILLER_34_701 VPWR VGND sg13g2_fill_2
XFILLER_33_200 VPWR VGND sg13g2_fill_2
X_4820_ VGND VPWR _1763_ _1764_ _1766_ _1758_ sg13g2_a21oi_1
XFILLER_22_929 VPWR VGND sg13g2_decap_8
X_4751_ _1693_ VPWR _1698_ VGND _1694_ _1696_ sg13g2_o21ai_1
XFILLER_21_439 VPWR VGND sg13g2_fill_2
XFILLER_30_951 VPWR VGND sg13g2_decap_8
X_3702_ VGND VPWR net578 _0861_ _0863_ _0862_ sg13g2_a21oi_1
X_4682_ _1630_ net756 net737 net762 net732 VPWR VGND sg13g2_a22oi_1
X_3633_ net576 VPWR _0800_ VGND _0798_ _0799_ sg13g2_o21ai_1
X_3564_ net584 _0624_ _0735_ VPWR VGND sg13g2_nor2_1
X_5303_ net94 VGND VPWR net377 ppwm_i.u_ppwm.data_o clknet_leaf_15_clk sg13g2_dfrbpq_1
X_3495_ _0657_ VPWR _0669_ VGND _0619_ _0658_ sg13g2_o21ai_1
X_5234_ net465 net626 _2141_ VPWR VGND sg13g2_nor2_1
X_5165_ _2101_ net1074 net777 net622 net1054 VPWR VGND sg13g2_a22oi_1
XFILLER_25_1002 VPWR VGND sg13g2_decap_8
X_4116_ falu_i.falutop.div_inst.acc\[1\] falu_i.falutop.div_inst.b1\[1\] _1118_ VPWR
+ VGND sg13g2_xor2_1
X_5096_ _2033_ _2020_ _2036_ VPWR VGND sg13g2_xor2_1
X_4047_ _1070_ _1069_ net985 _1068_ _1059_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_572 VPWR VGND sg13g2_fill_2
XFILLER_25_756 VPWR VGND sg13g2_fill_2
XFILLER_13_929 VPWR VGND sg13g2_decap_8
X_4949_ VPWR _1892_ _1891_ VGND sg13g2_inv_1
X_5510__245 VPWR VGND net245 sg13g2_tiehi
XFILLER_21_973 VPWR VGND sg13g2_decap_8
XFILLER_32_1017 VPWR VGND sg13g2_decap_8
XFILLER_32_1028 VPWR VGND sg13g2_fill_1
XFILLER_4_605 VPWR VGND sg13g2_decap_8
X_5252__191 VPWR VGND net191 sg13g2_tiehi
XFILLER_3_115 VPWR VGND sg13g2_fill_1
XFILLER_3_159 VPWR VGND sg13g2_fill_1
XFILLER_0_855 VPWR VGND sg13g2_decap_8
XFILLER_16_723 VPWR VGND sg13g2_decap_8
XFILLER_16_756 VPWR VGND sg13g2_fill_2
XFILLER_16_778 VPWR VGND sg13g2_decap_4
XFILLER_12_951 VPWR VGND sg13g2_decap_8
XFILLER_30_258 VPWR VGND sg13g2_fill_1
XFILLER_8_944 VPWR VGND sg13g2_decap_8
XFILLER_7_432 VPWR VGND sg13g2_fill_2
X_5571__56 VPWR VGND net56 sg13g2_tiehi
X_3280_ ppwm_i.u_ppwm.u_pwm.counter\[2\] _2286_ _0463_ VPWR VGND sg13g2_nor2_1
XFILLER_0_84 VPWR VGND sg13g2_decap_4
XFILLER_34_520 VPWR VGND sg13g2_fill_1
XFILLER_34_542 VPWR VGND sg13g2_fill_2
X_4803_ _1749_ _1699_ _1702_ VPWR VGND sg13g2_nand2_1
X_2995_ _2349_ net698 ppwm_i.u_ppwm.u_mem.memory\[58\] net703 ppwm_i.u_ppwm.u_mem.memory\[79\]
+ VPWR VGND sg13g2_a22oi_1
X_4734_ _1636_ VPWR _1681_ VGND _1550_ _1637_ sg13g2_o21ai_1
XFILLER_30_781 VPWR VGND sg13g2_fill_1
X_4665_ _1216_ _1314_ _1613_ VPWR VGND sg13g2_nor2_1
X_3616_ _0784_ _0782_ _0783_ VPWR VGND sg13g2_nand2b_1
X_4596_ _1480_ _1544_ _1545_ VPWR VGND sg13g2_nor2b_1
X_3547_ _0718_ VPWR _0719_ VGND _2244_ net599 sg13g2_o21ai_1
X_5544__363 VPWR VGND net363 sg13g2_tiehi
XFILLER_0_129 VPWR VGND sg13g2_decap_4
X_3478_ net609 _0633_ _0653_ VPWR VGND sg13g2_nor2b_1
X_5217_ _2128_ net388 net622 VPWR VGND sg13g2_nand2_1
XFILLER_28_14 VPWR VGND sg13g2_decap_8
XFILLER_29_303 VPWR VGND sg13g2_decap_4
X_5148_ net774 VPWR _2086_ VGND falu_i.falutop.div_inst.rem\[6\] _2047_ sg13g2_o21ai_1
X_5079_ _1997_ _1939_ _1996_ _2019_ VPWR VGND sg13g2_a21o_1
XFILLER_28_69 VPWR VGND sg13g2_fill_1
XFILLER_29_358 VPWR VGND sg13g2_decap_4
XFILLER_44_306 VPWR VGND sg13g2_fill_2
XFILLER_44_79 VPWR VGND sg13g2_fill_2
XFILLER_12_236 VPWR VGND sg13g2_decap_8
XFILLER_5_958 VPWR VGND sg13g2_decap_8
XFILLER_5_29 VPWR VGND sg13g2_fill_1
XFILLER_4_457 VPWR VGND sg13g2_decap_8
XFILLER_0_685 VPWR VGND sg13g2_decap_8
XFILLER_47_188 VPWR VGND sg13g2_fill_1
X_5376__300 VPWR VGND net300 sg13g2_tiehi
XFILLER_29_881 VPWR VGND sg13g2_fill_2
XFILLER_43_350 VPWR VGND sg13g2_fill_1
XFILLER_16_553 VPWR VGND sg13g2_decap_8
XFILLER_15_1001 VPWR VGND sg13g2_decap_8
XFILLER_34_90 VPWR VGND sg13g2_decap_4
XFILLER_8_741 VPWR VGND sg13g2_fill_2
XFILLER_12_792 VPWR VGND sg13g2_fill_1
XFILLER_7_284 VPWR VGND sg13g2_fill_2
X_4450_ _1370_ _1391_ _1360_ _1402_ VPWR VGND _1401_ sg13g2_nand4_1
Xhold207 _0239_ VPWR VGND net859 sg13g2_dlygate4sd3_1
X_3401_ VGND VPWR ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] _2261_ _0579_ _0578_ sg13g2_a21oi_1
X_4381_ VGND VPWR _2297_ net710 _1334_ net722 sg13g2_a21oi_1
Xhold229 falu_i.falutop.i2c_inst.data_in\[4\] VPWR VGND net881 sg13g2_dlygate4sd3_1
Xhold218 _0233_ VPWR VGND net870 sg13g2_dlygate4sd3_1
X_3332_ net1162 _0506_ _0511_ VPWR VGND sg13g2_nor2_1
Xfanout709 _2256_ net709 VPWR VGND sg13g2_buf_1
X_3263_ _2262_ _0449_ _0451_ VPWR VGND sg13g2_and2_1
XFILLER_39_634 VPWR VGND sg13g2_fill_2
X_5002_ net711 net766 net761 net755 _1944_ VPWR VGND sg13g2_and4_1
X_3194_ _0036_ net809 _0404_ net1050 VPWR VGND sg13g2_and3_1
XFILLER_22_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_188 VPWR VGND sg13g2_decap_8
XFILLER_27_829 VPWR VGND sg13g2_fill_1
X_5574__367 VPWR VGND net367 sg13g2_tiehi
Xclkbuf_3_5__f_clk clknet_0_clk clknet_3_5__leaf_clk VPWR VGND sg13g2_buf_8
X_2978_ VGND VPWR _2166_ net694 _2332_ net709 sg13g2_a21oi_1
X_4717_ _1664_ _1309_ _1662_ VPWR VGND sg13g2_nand2_1
X_4648_ _1533_ _1594_ _1530_ _1596_ VPWR VGND sg13g2_nand3_1
X_4579_ _1528_ net740 net710 VPWR VGND sg13g2_nand2_1
XFILLER_2_939 VPWR VGND sg13g2_decap_8
X_5299__99 VPWR VGND net99 sg13g2_tiehi
X_5310__81 VPWR VGND net81 sg13g2_tiehi
XFILLER_38_1023 VPWR VGND sg13g2_decap_4
XFILLER_13_501 VPWR VGND sg13g2_decap_4
XFILLER_26_895 VPWR VGND sg13g2_decap_8
XFILLER_9_516 VPWR VGND sg13g2_fill_1
XFILLER_40_386 VPWR VGND sg13g2_fill_2
XFILLER_5_755 VPWR VGND sg13g2_fill_2
XFILLER_4_221 VPWR VGND sg13g2_fill_1
XFILLER_20_70 VPWR VGND sg13g2_fill_2
XFILLER_45_1027 VPWR VGND sg13g2_fill_2
XFILLER_49_943 VPWR VGND sg13g2_decap_8
XFILLER_1_994 VPWR VGND sg13g2_decap_8
X_5301__92 VPWR VGND net92 sg13g2_tiehi
Xhold90 _0208_ VPWR VGND net462 sg13g2_dlygate4sd3_1
XFILLER_35_147 VPWR VGND sg13g2_fill_2
X_3950_ VGND VPWR _2168_ net677 _0194_ _1003_ sg13g2_a21oi_1
XFILLER_17_862 VPWR VGND sg13g2_decap_8
X_2901_ _2255_ net419 VPWR VGND sg13g2_inv_2
XFILLER_32_810 VPWR VGND sg13g2_fill_2
X_3881_ net840 VPWR _0969_ VGND ppwm_i.u_ppwm.u_mem.memory\[60\] net677 sg13g2_o21ai_1
XFILLER_31_320 VPWR VGND sg13g2_fill_1
XFILLER_32_854 VPWR VGND sg13g2_fill_2
X_2832_ VPWR _2186_ net463 VGND sg13g2_inv_1
X_5551_ net243 VGND VPWR net1030 falu_i.falutop.i2c_inst.result\[15\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_4502_ VGND VPWR _2296_ _1292_ _1453_ _1288_ sg13g2_a21oi_1
X_5482_ net321 VGND VPWR net895 falu_i.falutop.data_in\[13\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4433_ _1266_ _1235_ _1385_ VPWR VGND sg13g2_xor2_1
X_4364_ _1259_ _1279_ _1317_ VPWR VGND sg13g2_nor2_2
X_3315_ _0495_ net788 net701 VPWR VGND sg13g2_xnor2_1
X_4295_ _1248_ net632 _1246_ VPWR VGND sg13g2_xnor2_1
X_3246_ net1139 _0439_ _0440_ VPWR VGND sg13g2_and2_1
X_3177_ net813 VPWR _0394_ VGND ppwm_i.u_ppwm.pwm_value\[7\] net682 sg13g2_o21ai_1
X_5535__104 VPWR VGND net104 sg13g2_tiehi
XFILLER_41_128 VPWR VGND sg13g2_fill_1
XFILLER_23_821 VPWR VGND sg13g2_decap_8
XFILLER_25_48 VPWR VGND sg13g2_fill_1
XFILLER_23_898 VPWR VGND sg13g2_decap_8
XFILLER_10_537 VPWR VGND sg13g2_fill_2
XFILLER_2_703 VPWR VGND sg13g2_decap_8
XFILLER_2_747 VPWR VGND sg13g2_decap_4
XFILLER_46_902 VPWR VGND sg13g2_decap_8
XFILLER_46_979 VPWR VGND sg13g2_decap_8
XFILLER_26_681 VPWR VGND sg13g2_fill_1
XFILLER_13_342 VPWR VGND sg13g2_decap_4
XFILLER_14_887 VPWR VGND sg13g2_decap_8
X_3100_ VGND VPWR net800 net1002 _0005_ _2448_ sg13g2_a21oi_1
XFILLER_1_791 VPWR VGND sg13g2_decap_8
X_4080_ _1084_ _1082_ _1083_ _1081_ _1080_ VPWR VGND sg13g2_a22oi_1
XFILLER_49_784 VPWR VGND sg13g2_decap_4
XFILLER_37_902 VPWR VGND sg13g2_fill_2
X_3031_ VGND VPWR _2221_ net692 _2385_ net788 sg13g2_a21oi_1
XFILLER_37_957 VPWR VGND sg13g2_decap_8
XFILLER_24_607 VPWR VGND sg13g2_decap_4
X_4982_ net616 VPWR _1925_ VGND net739 net563 sg13g2_o21ai_1
XFILLER_16_191 VPWR VGND sg13g2_fill_2
X_3933_ net838 VPWR _0995_ VGND net544 net675 sg13g2_o21ai_1
X_3864_ VGND VPWR _2199_ net665 _0151_ _0960_ sg13g2_a21oi_1
X_2815_ VPWR _2169_ net867 VGND sg13g2_inv_1
XFILLER_20_846 VPWR VGND sg13g2_decap_8
X_5565__108 VPWR VGND net108 sg13g2_tiehi
X_3795_ net827 VPWR _0926_ VGND net447 net659 sg13g2_o21ai_1
X_5534_ net112 VGND VPWR net486 falu_i.falutop.div_inst.acc\[7\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_1
X_5465_ net361 VGND VPWR _0224_ falu_i.falutop.i2c_inst.counter\[2\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_4416_ VGND VPWR net707 net587 _1368_ _1367_ sg13g2_a21oi_1
X_5396_ net260 VGND VPWR _0155_ ppwm_i.u_ppwm.u_mem.memory\[55\] clknet_leaf_26_clk
+ sg13g2_dfrbpq_2
XFILLER_28_1022 VPWR VGND sg13g2_decap_8
X_5506__261 VPWR VGND net261 sg13g2_tiehi
X_4347_ net730 net735 net587 _1300_ VPWR VGND sg13g2_mux2_1
X_4278_ falu_i.falutop.alu_data_in\[9\] net767 _1231_ VPWR VGND sg13g2_nor2_2
XFILLER_28_924 VPWR VGND sg13g2_decap_8
X_3229_ _2271_ _0427_ _0429_ VPWR VGND sg13g2_and2_1
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_36_14 VPWR VGND sg13g2_decap_4
XFILLER_15_618 VPWR VGND sg13g2_decap_8
XFILLER_36_990 VPWR VGND sg13g2_decap_8
XFILLER_42_448 VPWR VGND sg13g2_decap_8
XFILLER_23_651 VPWR VGND sg13g2_decap_8
XFILLER_10_301 VPWR VGND sg13g2_fill_1
XFILLER_22_161 VPWR VGND sg13g2_decap_4
XFILLER_23_673 VPWR VGND sg13g2_decap_4
XFILLER_35_1026 VPWR VGND sg13g2_fill_2
XFILLER_11_846 VPWR VGND sg13g2_decap_8
XFILLER_7_839 VPWR VGND sg13g2_decap_8
Xhold390 _0302_ VPWR VGND net1042 sg13g2_dlygate4sd3_1
XFILLER_42_1008 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_decap_4
XFILLER_18_434 VPWR VGND sg13g2_fill_2
XFILLER_19_968 VPWR VGND sg13g2_decap_8
XFILLER_13_150 VPWR VGND sg13g2_fill_1
XFILLER_14_673 VPWR VGND sg13g2_decap_4
X_3580_ _0746_ _0749_ _0750_ VPWR VGND sg13g2_and2_1
XFILLER_6_850 VPWR VGND sg13g2_decap_8
XFILLER_5_382 VPWR VGND sg13g2_decap_4
X_5250_ net195 VGND VPWR _0012_ falu_i.falutop.i2c_inst.data_in\[8\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_1
X_5384__284 VPWR VGND net284 sg13g2_tiehi
X_4201_ VGND VPWR net633 _1171_ _0276_ _1172_ sg13g2_a21oi_1
X_5181_ net1123 net618 _2107_ VPWR VGND sg13g2_nor2_1
X_4132_ VPWR _0246_ net911 VGND sg13g2_inv_1
XFILLER_37_710 VPWR VGND sg13g2_decap_4
X_4063_ net881 falu_i.falutop.data_in\[4\] net685 _0232_ VPWR VGND sg13g2_mux2_1
X_3014_ _2368_ net688 ppwm_i.u_ppwm.u_mem.memory\[13\] net700 ppwm_i.u_ppwm.u_mem.memory\[27\]
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_765 VPWR VGND sg13g2_fill_2
XFILLER_36_253 VPWR VGND sg13g2_fill_1
XFILLER_36_286 VPWR VGND sg13g2_decap_4
X_4965_ net764 net755 net711 _1908_ VPWR VGND sg13g2_nand3_1
XFILLER_24_459 VPWR VGND sg13g2_decap_8
X_3916_ VGND VPWR _2180_ net669 _0177_ _0986_ sg13g2_a21oi_1
XFILLER_33_960 VPWR VGND sg13g2_decap_8
X_4896_ net815 VPWR _1840_ VGND net1064 net627 sg13g2_o21ai_1
X_3847_ net830 VPWR _0952_ VGND net860 net643 sg13g2_o21ai_1
XFILLER_20_698 VPWR VGND sg13g2_fill_2
X_3778_ VGND VPWR _2229_ net644 _0108_ _0917_ sg13g2_a21oi_1
X_5517_ net217 VGND VPWR _0276_ falu_i.falutop.div_inst.rem\[4\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_5448_ net98 VGND VPWR _0207_ ppwm_i.u_ppwm.u_mem.memory\[107\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
X_5379_ net294 VGND VPWR net423 ppwm_i.u_ppwm.u_mem.memory\[38\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
XFILLER_16_916 VPWR VGND sg13g2_decap_8
XFILLER_42_212 VPWR VGND sg13g2_decap_4
XFILLER_28_798 VPWR VGND sg13g2_fill_1
XFILLER_3_875 VPWR VGND sg13g2_decap_8
XFILLER_2_385 VPWR VGND sg13g2_fill_1
XFILLER_26_8 VPWR VGND sg13g2_fill_1
XFILLER_19_721 VPWR VGND sg13g2_fill_2
XFILLER_46_551 VPWR VGND sg13g2_fill_2
XFILLER_46_595 VPWR VGND sg13g2_decap_8
XFILLER_46_584 VPWR VGND sg13g2_fill_1
XFILLER_46_573 VPWR VGND sg13g2_fill_2
XFILLER_34_713 VPWR VGND sg13g2_fill_2
XFILLER_22_908 VPWR VGND sg13g2_decap_8
X_4750_ _1693_ _1694_ _1696_ _1697_ VPWR VGND sg13g2_or3_1
XFILLER_30_930 VPWR VGND sg13g2_decap_8
XFILLER_33_289 VPWR VGND sg13g2_fill_1
X_3701_ _0862_ _0740_ _0813_ VPWR VGND sg13g2_nand2_1
X_4681_ net738 net763 net732 _1629_ VPWR VGND net756 sg13g2_nand4_1
X_3632_ _0799_ ppwm_i.u_ppwm.pwm_value\[9\] net603 VPWR VGND sg13g2_xnor2_1
X_5302_ net90 VGND VPWR net1032 ppwm_i.u_ppwm.global_counter\[19\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
X_3563_ _0630_ _0694_ _0734_ VPWR VGND sg13g2_nor2_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_3494_ _0668_ _2250_ net600 VPWR VGND sg13g2_xnor2_1
X_5233_ _2092_ net775 _2140_ VPWR VGND sg13g2_nor2b_1
X_5164_ net1073 net622 _2099_ _2100_ VPWR VGND sg13g2_nor3_1
X_4115_ falu_i.falutop.div_inst.acc\[0\] falu_i.falutop.div_inst.b1\[0\] _1117_ VPWR
+ VGND sg13g2_nor2b_1
X_5095_ _2035_ _2020_ _2033_ VPWR VGND sg13g2_nand2_1
X_4046_ _1059_ VPWR _1069_ VGND _2440_ _1057_ sg13g2_o21ai_1
XFILLER_24_201 VPWR VGND sg13g2_decap_8
XFILLER_25_735 VPWR VGND sg13g2_decap_8
XFILLER_13_908 VPWR VGND sg13g2_decap_8
X_4948_ _1849_ VPWR _1891_ VGND _1795_ _1850_ sg13g2_o21ai_1
X_4879_ _1824_ _1790_ _1823_ VPWR VGND sg13g2_nand2_1
XFILLER_21_952 VPWR VGND sg13g2_decap_8
XFILLER_20_473 VPWR VGND sg13g2_fill_2
XFILLER_0_834 VPWR VGND sg13g2_decap_8
XFILLER_28_540 VPWR VGND sg13g2_decap_4
XFILLER_15_245 VPWR VGND sg13g2_decap_4
XFILLER_15_256 VPWR VGND sg13g2_fill_1
XFILLER_12_930 VPWR VGND sg13g2_decap_8
XFILLER_30_237 VPWR VGND sg13g2_fill_2
XFILLER_8_923 VPWR VGND sg13g2_decap_8
XFILLER_17_4 VPWR VGND sg13g2_fill_2
XFILLER_0_1016 VPWR VGND sg13g2_decap_8
XFILLER_0_1027 VPWR VGND sg13g2_fill_2
XFILLER_19_573 VPWR VGND sg13g2_decap_4
XFILLER_46_392 VPWR VGND sg13g2_fill_2
XFILLER_34_565 VPWR VGND sg13g2_fill_1
X_2994_ VGND VPWR ppwm_i.u_ppwm.u_mem.memory\[65\] net691 _2348_ net789 sg13g2_a21oi_1
X_4802_ _1748_ _1741_ _1746_ VPWR VGND sg13g2_xnor2_1
XFILLER_21_237 VPWR VGND sg13g2_fill_1
X_4733_ _1680_ _1638_ _1563_ VPWR VGND sg13g2_nand2b_1
X_4664_ _1612_ _1218_ _1611_ VPWR VGND sg13g2_xnor2_1
X_3615_ _0783_ _2244_ net603 VPWR VGND sg13g2_xnor2_1
X_4595_ _1542_ _1541_ _1544_ VPWR VGND sg13g2_xor2_1
X_3546_ _0718_ net782 net599 VPWR VGND sg13g2_nand2_1
X_5216_ falu_i.falutop.data_in\[8\] net906 net622 _0336_ VPWR VGND sg13g2_mux2_1
X_5427__184 VPWR VGND net184 sg13g2_tiehi
X_3477_ net584 net574 _0651_ _0652_ VPWR VGND sg13g2_nor3_1
X_5147_ _1590_ VPWR _2085_ VGND _2083_ _2084_ sg13g2_o21ai_1
X_5078_ _2017_ _2018_ _0307_ VPWR VGND sg13g2_nor2_1
XFILLER_38_871 VPWR VGND sg13g2_fill_2
X_4029_ _1054_ _1055_ _0221_ VPWR VGND sg13g2_nor2_1
XFILLER_37_381 VPWR VGND sg13g2_fill_2
XFILLER_9_709 VPWR VGND sg13g2_decap_4
X_5434__155 VPWR VGND net155 sg13g2_tiehi
X_5538__76 VPWR VGND net76 sg13g2_tiehi
XFILLER_5_937 VPWR VGND sg13g2_decap_8
X_5459__50 VPWR VGND net50 sg13g2_tiehi
X_5441__126 VPWR VGND net126 sg13g2_tiehi
XFILLER_35_307 VPWR VGND sg13g2_decap_4
XFILLER_16_565 VPWR VGND sg13g2_fill_1
XFILLER_12_771 VPWR VGND sg13g2_decap_4
XFILLER_7_241 VPWR VGND sg13g2_decap_4
Xhold208 ppwm_i.u_ppwm.u_mem.memory\[44\] VPWR VGND net860 sg13g2_dlygate4sd3_1
X_3400_ VPWR VGND _2238_ _0577_ ppwm_i.u_ppwm.global_counter\[15\] _2237_ _0578_ ppwm_i.u_ppwm.global_counter\[16\]
+ sg13g2_a221oi_1
Xhold219 falu_i.falutop.i2c_inst.data_in\[7\] VPWR VGND net871 sg13g2_dlygate4sd3_1
X_4380_ _1285_ _1332_ _1333_ VPWR VGND sg13g2_and2_1
X_3331_ _0509_ _0508_ _0510_ VPWR VGND sg13g2_xor2_1
XFILLER_4_992 VPWR VGND sg13g2_decap_8
X_3262_ net975 _0450_ _0059_ VPWR VGND sg13g2_nor2_1
X_5001_ _1943_ _1897_ _1942_ VPWR VGND sg13g2_xnor2_1
XFILLER_22_1006 VPWR VGND sg13g2_decap_8
X_3193_ _0405_ net1049 _0402_ VPWR VGND sg13g2_nand2_1
XFILLER_26_307 VPWR VGND sg13g2_fill_2
XFILLER_34_340 VPWR VGND sg13g2_fill_1
X_2977_ _2331_ _2171_ net690 VPWR VGND sg13g2_nand2_1
X_4716_ VGND VPWR _1602_ _1605_ _1663_ _1661_ sg13g2_a21oi_1
X_4647_ _1533_ _1530_ _1594_ _1595_ VPWR VGND sg13g2_a21o_2
XFILLER_30_16 VPWR VGND sg13g2_fill_1
X_4578_ _1527_ net731 net721 VPWR VGND sg13g2_nand2_1
XFILLER_2_918 VPWR VGND sg13g2_decap_8
X_3529_ VPWR VGND _0622_ _0698_ _0701_ net571 _0702_ _0648_ sg13g2_a221oi_1
XFILLER_29_145 VPWR VGND sg13g2_fill_2
XFILLER_26_830 VPWR VGND sg13g2_decap_8
XFILLER_38_1002 VPWR VGND sg13g2_decap_8
XFILLER_26_874 VPWR VGND sg13g2_decap_8
XFILLER_40_343 VPWR VGND sg13g2_fill_1
XFILLER_40_332 VPWR VGND sg13g2_decap_8
XFILLER_5_745 VPWR VGND sg13g2_fill_2
XFILLER_4_211 VPWR VGND sg13g2_fill_1
XFILLER_45_1006 VPWR VGND sg13g2_decap_8
XFILLER_49_922 VPWR VGND sg13g2_decap_8
XFILLER_1_973 VPWR VGND sg13g2_decap_8
X_5343__366 VPWR VGND net366 sg13g2_tiehi
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_49_999 VPWR VGND sg13g2_decap_8
XFILLER_48_465 VPWR VGND sg13g2_fill_1
Xhold91 ppwm_i.u_ppwm.u_mem.memory\[70\] VPWR VGND net463 sg13g2_dlygate4sd3_1
Xhold80 falu_i.falutop.div_inst.a\[4\] VPWR VGND net452 sg13g2_dlygate4sd3_1
XFILLER_17_841 VPWR VGND sg13g2_decap_8
XFILLER_35_115 VPWR VGND sg13g2_decap_4
XFILLER_36_638 VPWR VGND sg13g2_fill_1
XFILLER_44_671 VPWR VGND sg13g2_fill_1
X_2900_ net786 _2254_ VPWR VGND sg13g2_inv_4
X_3880_ VGND VPWR _2193_ net676 _0159_ _0968_ sg13g2_a21oi_1
XFILLER_43_192 VPWR VGND sg13g2_fill_1
XFILLER_16_395 VPWR VGND sg13g2_fill_1
XFILLER_31_332 VPWR VGND sg13g2_fill_1
X_2831_ VPWR _2185_ net415 VGND sg13g2_inv_1
XFILLER_31_365 VPWR VGND sg13g2_fill_1
X_5550_ net251 VGND VPWR net1072 falu_i.falutop.i2c_inst.result\[14\] clknet_leaf_42_clk
+ sg13g2_dfrbpq_1
X_5481_ net323 VGND VPWR net927 falu_i.falutop.data_in\[12\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4501_ _1452_ net587 net725 VPWR VGND sg13g2_nand2b_1
X_4432_ _1384_ _1234_ _1383_ VPWR VGND sg13g2_nand2_1
X_4363_ _1316_ _1315_ _1221_ VPWR VGND sg13g2_nand2b_1
X_4294_ VGND VPWR _1247_ _1245_ _1243_ sg13g2_or2_1
X_5540__60 VPWR VGND net60 sg13g2_tiehi
X_3314_ _0067_ _0492_ _0494_ VPWR VGND sg13g2_nand2_1
X_3245_ net795 net554 _0439_ _0053_ VPWR VGND sg13g2_nor3_1
XFILLER_6_1011 VPWR VGND sg13g2_decap_8
X_3176_ VGND VPWR _2282_ net682 _0030_ _0393_ sg13g2_a21oi_1
XFILLER_39_465 VPWR VGND sg13g2_fill_1
XFILLER_39_454 VPWR VGND sg13g2_decap_8
X_5394__264 VPWR VGND net264 sg13g2_tiehi
XFILLER_23_800 VPWR VGND sg13g2_decap_8
XFILLER_25_16 VPWR VGND sg13g2_fill_1
XFILLER_41_118 VPWR VGND sg13g2_fill_1
XFILLER_23_877 VPWR VGND sg13g2_decap_8
X_5249__197 VPWR VGND net197 sg13g2_tiehi
XFILLER_46_958 VPWR VGND sg13g2_decap_8
XFILLER_17_148 VPWR VGND sg13g2_decap_4
X_5553__227 VPWR VGND net227 sg13g2_tiehi
XFILLER_33_619 VPWR VGND sg13g2_decap_8
XFILLER_14_866 VPWR VGND sg13g2_decap_8
XFILLER_41_696 VPWR VGND sg13g2_fill_2
XFILLER_5_520 VPWR VGND sg13g2_fill_1
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_5_597 VPWR VGND sg13g2_fill_2
XFILLER_49_741 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_decap_8
X_3030_ VPWR VGND _2202_ _2382_ net692 _2197_ _2384_ net700 sg13g2_a221oi_1
XFILLER_48_295 VPWR VGND sg13g2_fill_1
XFILLER_37_936 VPWR VGND sg13g2_decap_8
XFILLER_36_457 VPWR VGND sg13g2_decap_8
XFILLER_36_479 VPWR VGND sg13g2_fill_1
X_4981_ net765 net563 _1924_ VPWR VGND sg13g2_nor2b_1
Xclkbuf_leaf_43_clk clknet_3_0__leaf_clk clknet_leaf_43_clk VPWR VGND sg13g2_buf_8
XFILLER_32_630 VPWR VGND sg13g2_decap_8
X_3932_ VGND VPWR _2174_ net650 _0185_ _0994_ sg13g2_a21oi_1
X_3863_ net830 VPWR _0960_ VGND ppwm_i.u_ppwm.u_mem.memory\[51\] net665 sg13g2_o21ai_1
XFILLER_20_825 VPWR VGND sg13g2_decap_8
XFILLER_32_663 VPWR VGND sg13g2_decap_8
X_2814_ VPWR _2168_ net556 VGND sg13g2_inv_1
X_5533_ net120 VGND VPWR net932 falu_i.falutop.div_inst.acc\[6\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_9_881 VPWR VGND sg13g2_decap_8
X_3794_ VGND VPWR _2223_ net659 _0116_ _0925_ sg13g2_a21oi_1
X_5464_ net365 VGND VPWR _0223_ falu_i.falutop.i2c_inst.counter\[1\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_5395_ net262 VGND VPWR _0154_ ppwm_i.u_ppwm.u_mem.memory\[54\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4415_ net736 net587 _1367_ VPWR VGND sg13g2_nor2_1
XFILLER_28_1001 VPWR VGND sg13g2_decap_8
X_4346_ _1289_ _1298_ _1299_ VPWR VGND sg13g2_nor2_2
X_4277_ _1230_ _1228_ VPWR VGND _1226_ sg13g2_nand2b_2
XFILLER_39_240 VPWR VGND sg13g2_decap_4
XFILLER_28_903 VPWR VGND sg13g2_decap_8
X_3228_ VGND VPWR _2272_ _0425_ _0047_ _0428_ sg13g2_a21oi_1
XFILLER_39_284 VPWR VGND sg13g2_fill_2
X_3159_ net807 net373 _0023_ VPWR VGND sg13g2_and2_1
XFILLER_42_438 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_34_clk clknet_3_5__leaf_clk clknet_leaf_34_clk VPWR VGND sg13g2_buf_8
X_5513__233 VPWR VGND net233 sg13g2_tiehi
XFILLER_22_140 VPWR VGND sg13g2_decap_8
XFILLER_23_685 VPWR VGND sg13g2_decap_8
XFILLER_35_1005 VPWR VGND sg13g2_decap_8
XFILLER_7_807 VPWR VGND sg13g2_fill_2
XFILLER_10_335 VPWR VGND sg13g2_fill_1
Xhold380 _0064_ VPWR VGND net1032 sg13g2_dlygate4sd3_1
XFILLER_2_578 VPWR VGND sg13g2_decap_4
Xhold391 falu_i.falutop.i2c_inst.counter\[0\] VPWR VGND net1043 sg13g2_dlygate4sd3_1
X_5262__172 VPWR VGND net172 sg13g2_tiehi
XFILLER_19_947 VPWR VGND sg13g2_decap_8
XFILLER_27_980 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_25_clk clknet_3_6__leaf_clk clknet_leaf_25_clk VPWR VGND sg13g2_buf_8
XFILLER_14_641 VPWR VGND sg13g2_fill_1
XFILLER_14_652 VPWR VGND sg13g2_decap_8
XFILLER_42_994 VPWR VGND sg13g2_decap_8
XFILLER_9_133 VPWR VGND sg13g2_fill_2
XFILLER_14_696 VPWR VGND sg13g2_fill_2
X_5338__30 VPWR VGND net30 sg13g2_tiehi
XFILLER_10_880 VPWR VGND sg13g2_decap_8
X_4200_ net803 VPWR _1172_ VGND net1124 net635 sg13g2_o21ai_1
X_5180_ net1158 net743 net618 _0321_ VPWR VGND sg13g2_mux2_1
X_4131_ _1133_ net567 _1097_ net607 net910 VPWR VGND sg13g2_a22oi_1
XFILLER_3_74 VPWR VGND sg13g2_fill_1
XFILLER_49_560 VPWR VGND sg13g2_decap_4
X_4062_ net992 falu_i.falutop.data_in\[3\] net685 _0231_ VPWR VGND sg13g2_mux2_1
X_3013_ _2367_ _2364_ _2366_ _2363_ _2362_ VPWR VGND sg13g2_a22oi_1
XFILLER_36_232 VPWR VGND sg13g2_decap_8
XFILLER_18_991 VPWR VGND sg13g2_decap_8
XFILLER_25_939 VPWR VGND sg13g2_decap_8
XFILLER_36_276 VPWR VGND sg13g2_fill_1
Xclkbuf_leaf_16_clk clknet_3_2__leaf_clk clknet_leaf_16_clk VPWR VGND sg13g2_buf_8
X_4964_ net712 VPWR _1907_ VGND net761 net755 sg13g2_o21ai_1
X_3915_ net834 VPWR _0986_ VGND ppwm_i.u_ppwm.u_mem.memory\[77\] net669 sg13g2_o21ai_1
X_4895_ _1838_ _1839_ _0303_ VPWR VGND sg13g2_nor2_1
X_3846_ VGND VPWR _2205_ net665 _0142_ _0951_ sg13g2_a21oi_1
XFILLER_20_644 VPWR VGND sg13g2_decap_8
X_3777_ net830 VPWR _0917_ VGND ppwm_i.u_ppwm.u_mem.memory\[9\] net644 sg13g2_o21ai_1
X_5516_ net221 VGND VPWR _0275_ falu_i.falutop.div_inst.rem\[3\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_1
X_5447_ net102 VGND VPWR net446 ppwm_i.u_ppwm.u_mem.memory\[106\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_5378_ net296 VGND VPWR net425 ppwm_i.u_ppwm.u_mem.memory\[37\] clknet_leaf_21_clk
+ sg13g2_dfrbpq_1
X_4329_ _1282_ falu_i.falutop.alu_inst.op\[3\] _1280_ VPWR VGND sg13g2_nand2_2
XFILLER_47_508 VPWR VGND sg13g2_decap_4
XFILLER_47_14 VPWR VGND sg13g2_fill_1
XFILLER_43_725 VPWR VGND sg13g2_fill_1
XFILLER_42_235 VPWR VGND sg13g2_decap_8
XFILLER_11_622 VPWR VGND sg13g2_decap_8
XFILLER_7_648 VPWR VGND sg13g2_decap_8
XFILLER_6_114 VPWR VGND sg13g2_decap_8
XFILLER_7_659 VPWR VGND sg13g2_fill_2
X_5335__33 VPWR VGND net33 sg13g2_tiehi
XFILLER_5_0 VPWR VGND sg13g2_fill_1
XFILLER_3_854 VPWR VGND sg13g2_decap_8
XFILLER_19_700 VPWR VGND sg13g2_decap_4
Xfanout690 net691 net690 VPWR VGND sg13g2_buf_8
XFILLER_19_744 VPWR VGND sg13g2_fill_2
XFILLER_19_766 VPWR VGND sg13g2_decap_8
XFILLER_33_202 VPWR VGND sg13g2_fill_1
X_5494__291 VPWR VGND net291 sg13g2_tiehi
XFILLER_33_224 VPWR VGND sg13g2_decap_8
XFILLER_34_758 VPWR VGND sg13g2_decap_4
XFILLER_33_268 VPWR VGND sg13g2_fill_1
X_3700_ ppwm_i.u_ppwm.pwm_value\[5\] _0742_ net581 _0861_ VPWR VGND sg13g2_mux2_1
XFILLER_14_482 VPWR VGND sg13g2_fill_2
XFILLER_15_994 VPWR VGND sg13g2_decap_8
XFILLER_14_493 VPWR VGND sg13g2_decap_8
X_4680_ _1628_ _1557_ _1555_ VPWR VGND sg13g2_nand2b_1
X_3631_ VGND VPWR ppwm_i.u_ppwm.pwm_value\[8\] net603 _0798_ _0785_ sg13g2_a21oi_1
XFILLER_30_986 VPWR VGND sg13g2_decap_8
X_3562_ _0655_ _0714_ _0733_ VPWR VGND sg13g2_nor2_1
X_5301_ net92 VGND VPWR net1077 ppwm_i.u_ppwm.global_counter\[18\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
X_3493_ VGND VPWR _0656_ _0666_ _0073_ _0667_ sg13g2_a21oi_1
X_5232_ VGND VPWR net625 _2139_ _0340_ _2137_ sg13g2_a21oi_1
Xclkbuf_leaf_5_clk clknet_3_3__leaf_clk clknet_leaf_5_clk VPWR VGND sg13g2_buf_8
X_5163_ _2099_ _2098_ falu_i.falutop.data_in\[5\] VPWR VGND sg13g2_nand2b_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_4114_ _1116_ falu_i.falutop.div_inst.acc\[1\] falu_i.falutop.div_inst.b1\[1\] VPWR
+ VGND sg13g2_nand2b_1
X_5094_ _2020_ _2033_ _2034_ VPWR VGND sg13g2_nor2_1
X_4045_ _1068_ _1051_ _1067_ VPWR VGND sg13g2_nand2_1
XFILLER_25_703 VPWR VGND sg13g2_fill_1
XFILLER_25_714 VPWR VGND sg13g2_decap_8
XFILLER_25_758 VPWR VGND sg13g2_fill_1
XFILLER_40_717 VPWR VGND sg13g2_fill_1
XFILLER_12_408 VPWR VGND sg13g2_decap_8
XFILLER_40_739 VPWR VGND sg13g2_fill_2
X_4947_ _1872_ VPWR _1890_ VGND _1842_ _1873_ sg13g2_o21ai_1
XFILLER_21_931 VPWR VGND sg13g2_decap_8
X_4878_ _1823_ _1799_ _1822_ VPWR VGND sg13g2_xnor2_1
XFILLER_32_290 VPWR VGND sg13g2_fill_1
X_3829_ net825 VPWR _0943_ VGND net897 net656 sg13g2_o21ai_1
XFILLER_3_106 VPWR VGND sg13g2_decap_8
XFILLER_0_813 VPWR VGND sg13g2_decap_8
XFILLER_28_563 VPWR VGND sg13g2_fill_2
XFILLER_15_213 VPWR VGND sg13g2_decap_8
XFILLER_8_902 VPWR VGND sg13g2_decap_8
XFILLER_12_986 VPWR VGND sg13g2_decap_8
XFILLER_8_979 VPWR VGND sg13g2_decap_8
XFILLER_7_434 VPWR VGND sg13g2_fill_1
XFILLER_48_1026 VPWR VGND sg13g2_fill_2
XFILLER_31_7 VPWR VGND sg13g2_fill_2
XFILLER_39_806 VPWR VGND sg13g2_fill_2
XFILLER_38_349 VPWR VGND sg13g2_fill_2
XFILLER_38_338 VPWR VGND sg13g2_decap_8
XFILLER_47_883 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_34_500 VPWR VGND sg13g2_decap_4
XFILLER_34_544 VPWR VGND sg13g2_fill_1
XFILLER_22_706 VPWR VGND sg13g2_fill_2
X_2993_ _2347_ ppwm_i.u_ppwm.u_mem.memory\[72\] net695 VPWR VGND sg13g2_nand2_1
X_4801_ _1747_ _1741_ _1746_ VPWR VGND sg13g2_nand2_1
XFILLER_21_216 VPWR VGND sg13g2_fill_1
XFILLER_22_728 VPWR VGND sg13g2_decap_8
X_5353__346 VPWR VGND net346 sg13g2_tiehi
XFILLER_9_51 VPWR VGND sg13g2_decap_8
XFILLER_9_62 VPWR VGND sg13g2_fill_2
X_4732_ _1678_ VPWR _1679_ VGND _1567_ _1640_ sg13g2_o21ai_1
X_4663_ _1236_ _1572_ _1611_ VPWR VGND sg13g2_nor2_1
X_3614_ _0782_ _0747_ _0780_ _0781_ VPWR VGND sg13g2_and3_2
X_4594_ _1541_ _1542_ _1543_ VPWR VGND sg13g2_and2_1
X_3545_ _0716_ VPWR _0717_ VGND net584 _0626_ sg13g2_o21ai_1
X_3476_ VGND VPWR _0650_ _0651_ net598 ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] sg13g2_a21oi_2
X_5215_ VGND VPWR net623 _2127_ _0335_ _2126_ sg13g2_a21oi_1
X_5146_ _1834_ VPWR _2084_ VGND _1240_ _1282_ sg13g2_o21ai_1
X_5077_ net815 VPWR _2018_ VGND net1018 net627 sg13g2_o21ai_1
X_4028_ net816 VPWR _1055_ VGND net459 _1053_ sg13g2_o21ai_1
XFILLER_12_205 VPWR VGND sg13g2_decap_4
XFILLER_40_558 VPWR VGND sg13g2_decap_4
XFILLER_40_547 VPWR VGND sg13g2_decap_4
XFILLER_21_761 VPWR VGND sg13g2_fill_1
XFILLER_5_916 VPWR VGND sg13g2_decap_8
XFILLER_4_426 VPWR VGND sg13g2_decap_8
XFILLER_47_113 VPWR VGND sg13g2_decap_8
XFILLER_47_179 VPWR VGND sg13g2_fill_2
XFILLER_16_533 VPWR VGND sg13g2_fill_2
XFILLER_18_82 VPWR VGND sg13g2_decap_8
XFILLER_28_393 VPWR VGND sg13g2_decap_4
X_5259__177 VPWR VGND net177 sg13g2_tiehi
XFILLER_16_588 VPWR VGND sg13g2_decap_8
XFILLER_31_536 VPWR VGND sg13g2_fill_2
XFILLER_8_710 VPWR VGND sg13g2_decap_8
Xhold209 falu_i.falutop.i2c_inst.data_in\[14\] VPWR VGND net861 sg13g2_dlygate4sd3_1
X_3330_ _0497_ VPWR _0509_ VGND _0496_ _0498_ sg13g2_o21ai_1
XFILLER_4_971 VPWR VGND sg13g2_decap_8
X_5000_ _1942_ _1936_ _1940_ VPWR VGND sg13g2_xnor2_1
X_3261_ _0450_ net812 _0449_ VPWR VGND sg13g2_nand2_1
XFILLER_39_636 VPWR VGND sg13g2_fill_1
XFILLER_38_102 VPWR VGND sg13g2_decap_8
X_3192_ VGND VPWR _0404_ _0402_ net1049 sg13g2_or2_1
XFILLER_35_886 VPWR VGND sg13g2_fill_1
X_5470__345 VPWR VGND net345 sg13g2_tiehi
X_2976_ VPWR _2330_ _2329_ VGND sg13g2_inv_1
X_4715_ _1605_ _1661_ _1602_ _1662_ VPWR VGND sg13g2_nand3_1
X_4646_ VGND VPWR _1594_ _1593_ _1592_ sg13g2_or2_1
X_4577_ _1520_ _1521_ _1526_ _0298_ VPWR VGND sg13g2_nor3_1
X_3528_ _0677_ _0700_ net610 _0701_ VPWR VGND sg13g2_mux2_1
X_3459_ _0634_ VPWR _0635_ VGND net611 _0631_ sg13g2_o21ai_1
X_5129_ net749 net563 _2068_ VPWR VGND sg13g2_nor2b_1
XFILLER_26_842 VPWR VGND sg13g2_fill_2
XFILLER_26_853 VPWR VGND sg13g2_decap_8
XFILLER_13_547 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_13_569 VPWR VGND sg13g2_fill_1
XFILLER_5_713 VPWR VGND sg13g2_decap_4
XFILLER_5_757 VPWR VGND sg13g2_fill_1
XFILLER_4_267 VPWR VGND sg13g2_fill_1
XFILLER_20_72 VPWR VGND sg13g2_fill_1
XFILLER_49_901 VPWR VGND sg13g2_decap_8
XFILLER_1_952 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_49_978 VPWR VGND sg13g2_decap_8
Xhold92 _0169_ VPWR VGND net464 sg13g2_dlygate4sd3_1
Xhold81 _0340_ VPWR VGND net453 sg13g2_dlygate4sd3_1
Xhold70 _0108_ VPWR VGND net442 sg13g2_dlygate4sd3_1
XFILLER_17_820 VPWR VGND sg13g2_decap_8
XFILLER_35_149 VPWR VGND sg13g2_fill_1
XFILLER_16_352 VPWR VGND sg13g2_fill_1
XFILLER_17_897 VPWR VGND sg13g2_decap_8
X_2830_ VPWR _2184_ net977 VGND sg13g2_inv_1
XFILLER_31_311 VPWR VGND sg13g2_decap_8
XFILLER_31_344 VPWR VGND sg13g2_decap_4
X_5272__152 VPWR VGND net152 sg13g2_tiehi
XFILLER_31_388 VPWR VGND sg13g2_fill_1
XFILLER_31_399 VPWR VGND sg13g2_fill_2
X_5480_ net325 VGND VPWR net859 falu_i.falutop.data_in\[11\] clknet_leaf_38_clk sg13g2_dfrbpq_2
X_4500_ VGND VPWR _1297_ _1363_ _1451_ _1299_ sg13g2_a21oi_1
X_4431_ net772 _1303_ _1383_ VPWR VGND sg13g2_and2_1
X_4362_ _1312_ _1314_ _1307_ _1315_ VPWR VGND sg13g2_nand3_1
X_4293_ _1243_ _1245_ _1246_ VPWR VGND sg13g2_nor2_2
X_3313_ _0494_ net791 _0493_ VPWR VGND sg13g2_nand2_1
X_3244_ _2267_ _2268_ _2269_ _0433_ _0439_ VPWR VGND sg13g2_nor4_1
XFILLER_39_433 VPWR VGND sg13g2_decap_4
XFILLER_39_422 VPWR VGND sg13g2_fill_1
X_3175_ net810 VPWR _0393_ VGND ppwm_i.u_ppwm.pwm_value\[6\] net682 sg13g2_o21ai_1
XFILLER_23_856 VPWR VGND sg13g2_decap_8
XFILLER_34_171 VPWR VGND sg13g2_fill_1
X_2959_ _2313_ net794 net791 VPWR VGND sg13g2_nand2b_1
X_4629_ _1578_ _1577_ _1576_ VPWR VGND sg13g2_nand2b_1
Xhold540 ppwm_i.u_ppwm.pc\[3\] VPWR VGND net1192 sg13g2_dlygate4sd3_1
XFILLER_2_716 VPWR VGND sg13g2_decap_4
XFILLER_45_403 VPWR VGND sg13g2_fill_1
XFILLER_18_617 VPWR VGND sg13g2_fill_2
XFILLER_46_937 VPWR VGND sg13g2_decap_8
XFILLER_14_845 VPWR VGND sg13g2_decap_8
XFILLER_41_675 VPWR VGND sg13g2_decap_8
XFILLER_13_355 VPWR VGND sg13g2_fill_2
XFILLER_12_1028 VPWR VGND sg13g2_fill_1
XFILLER_5_565 VPWR VGND sg13g2_decap_4
XFILLER_5_576 VPWR VGND sg13g2_fill_1
XFILLER_36_436 VPWR VGND sg13g2_decap_8
XFILLER_45_992 VPWR VGND sg13g2_decap_8
X_4980_ _1318_ _1921_ _1922_ _1923_ VPWR VGND sg13g2_nor3_2
XFILLER_23_119 VPWR VGND sg13g2_fill_2
XFILLER_16_182 VPWR VGND sg13g2_fill_1
X_3931_ net837 VPWR _0994_ VGND ppwm_i.u_ppwm.u_mem.memory\[86\] net650 sg13g2_o21ai_1
X_3862_ VGND VPWR _2200_ net645 _0150_ _0959_ sg13g2_a21oi_1
XFILLER_20_804 VPWR VGND sg13g2_decap_8
X_2813_ VPWR _2167_ net532 VGND sg13g2_inv_1
X_5532_ net128 VGND VPWR net550 falu_i.falutop.div_inst.acc\[5\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_9_860 VPWR VGND sg13g2_decap_8
X_3793_ net828 VPWR _0925_ VGND ppwm_i.u_ppwm.u_mem.memory\[16\] net659 sg13g2_o21ai_1
X_5463_ net369 VGND VPWR _0222_ falu_i.falutop.i2c_inst.counter\[0\] clknet_leaf_5_clk
+ sg13g2_dfrbpq_2
X_5394_ net264 VGND VPWR _0153_ ppwm_i.u_ppwm.u_mem.memory\[53\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_4414_ net725 net730 net587 _1366_ VPWR VGND sg13g2_mux2_1
X_4345_ falu_i.falutop.alu_inst.op\[0\] _2299_ falu_i.falutop.alu_inst.op\[1\] _1298_
+ VPWR VGND net771 sg13g2_nand4_1
X_4276_ _1226_ _1227_ _1229_ VPWR VGND sg13g2_nor2_2
X_3227_ _0428_ net812 _0427_ VPWR VGND sg13g2_nand2_1
XFILLER_39_274 VPWR VGND sg13g2_decap_4
X_3158_ VGND VPWR net801 _0382_ _0022_ _0383_ sg13g2_a21oi_1
XFILLER_28_959 VPWR VGND sg13g2_decap_8
XFILLER_43_907 VPWR VGND sg13g2_fill_2
XFILLER_15_609 VPWR VGND sg13g2_decap_4
XFILLER_27_447 VPWR VGND sg13g2_fill_1
X_3089_ _2439_ _2433_ _2438_ VPWR VGND sg13g2_nand2_2
XFILLER_35_1028 VPWR VGND sg13g2_fill_1
XFILLER_6_318 VPWR VGND sg13g2_decap_4
XFILLER_7_4 VPWR VGND sg13g2_decap_8
Xhold381 falu_i.falutop.i2c_inst.result\[8\] VPWR VGND net1033 sg13g2_dlygate4sd3_1
Xhold370 falu_i.falutop.i2c_inst.result\[0\] VPWR VGND net1022 sg13g2_dlygate4sd3_1
Xhold392 falu_i.falutop.i2c_inst.data_in\[18\] VPWR VGND net1044 sg13g2_dlygate4sd3_1
XFILLER_19_926 VPWR VGND sg13g2_decap_8
XFILLER_33_406 VPWR VGND sg13g2_fill_1
XFILLER_42_973 VPWR VGND sg13g2_decap_8
XFILLER_9_167 VPWR VGND sg13g2_fill_2
XFILLER_9_178 VPWR VGND sg13g2_fill_1
XFILLER_6_885 VPWR VGND sg13g2_decap_8
XFILLER_5_362 VPWR VGND sg13g2_fill_1
XFILLER_5_395 VPWR VGND sg13g2_fill_2
X_4130_ _1131_ VPWR _1132_ VGND falu_i.falutop.div_inst.b1\[7\] _2290_ sg13g2_o21ai_1
X_4061_ net972 falu_i.falutop.data_in\[2\] net685 _0230_ VPWR VGND sg13g2_mux2_1
X_3012_ VPWR VGND ppwm_i.u_ppwm.u_mem.memory\[76\] _2365_ net694 ppwm_i.u_ppwm.u_mem.memory\[62\]
+ _2366_ net697 sg13g2_a221oi_1
XFILLER_3_1015 VPWR VGND sg13g2_decap_8
XFILLER_18_970 VPWR VGND sg13g2_decap_8
XFILLER_25_918 VPWR VGND sg13g2_decap_8
X_4963_ _1906_ _1214_ _1905_ VPWR VGND sg13g2_xnor2_1
X_3914_ VGND VPWR _2181_ net670 _0176_ _0985_ sg13g2_a21oi_1
X_4894_ net815 VPWR _1839_ VGND net1033 net627 sg13g2_o21ai_1
XFILLER_20_612 VPWR VGND sg13g2_fill_1
XFILLER_33_995 VPWR VGND sg13g2_decap_8
X_3845_ net829 VPWR _0951_ VGND ppwm_i.u_ppwm.u_mem.memory\[42\] net665 sg13g2_o21ai_1
XFILLER_22_18 VPWR VGND sg13g2_decap_8
X_3776_ VGND VPWR _2229_ net662 _0107_ _0916_ sg13g2_a21oi_1
X_5515_ net225 VGND VPWR _0274_ falu_i.falutop.div_inst.rem\[2\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_5446_ net106 VGND VPWR net529 ppwm_i.u_ppwm.u_mem.memory\[105\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_1
X_5363__326 VPWR VGND net326 sg13g2_tiehi
X_5377_ net298 VGND VPWR _0136_ ppwm_i.u_ppwm.u_mem.memory\[36\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_4328_ net772 _2300_ _1279_ _1281_ VPWR VGND sg13g2_nor3_2
X_4259_ _1213_ _1182_ _1097_ net607 net879 VPWR VGND sg13g2_a22oi_1
XFILLER_27_200 VPWR VGND sg13g2_fill_2
XFILLER_28_723 VPWR VGND sg13g2_decap_8
XFILLER_15_417 VPWR VGND sg13g2_fill_2
X_5437__143 VPWR VGND net143 sg13g2_tiehi
XFILLER_15_439 VPWR VGND sg13g2_decap_4
XFILLER_24_984 VPWR VGND sg13g2_decap_8
XFILLER_7_627 VPWR VGND sg13g2_fill_2
X_5409__234 VPWR VGND net234 sg13g2_tiehi
XFILLER_3_833 VPWR VGND sg13g2_decap_8
X_5444__114 VPWR VGND net114 sg13g2_tiehi
Xfanout691 _2312_ net691 VPWR VGND sg13g2_buf_8
XFILLER_19_723 VPWR VGND sg13g2_fill_1
Xfanout680 net884 net680 VPWR VGND sg13g2_buf_8
XFILLER_18_211 VPWR VGND sg13g2_decap_8
XFILLER_18_222 VPWR VGND sg13g2_fill_2
XFILLER_34_715 VPWR VGND sg13g2_fill_1
XFILLER_15_973 VPWR VGND sg13g2_decap_8
XFILLER_18_1012 VPWR VGND sg13g2_decap_8
XFILLER_33_258 VPWR VGND sg13g2_decap_4
XFILLER_30_965 VPWR VGND sg13g2_decap_8
X_3630_ VPWR VGND _0797_ net799 _0786_ _2244_ _0080_ net573 sg13g2_a221oi_1
X_3561_ _0730_ _0731_ net575 _0732_ VPWR VGND sg13g2_nand3_1
X_5300_ net97 VGND VPWR net991 ppwm_i.u_ppwm.global_counter\[17\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_2
X_3492_ net821 VPWR _0667_ VGND net784 _0614_ sg13g2_o21ai_1
X_5231_ _2139_ falu_i.falutop.data_in\[12\] _2138_ VPWR VGND sg13g2_xnor2_1
X_5162_ falu_i.falutop.data_in\[4\] _2097_ _2098_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_1016 VPWR VGND sg13g2_decap_8
X_5093_ _2033_ _2023_ _2032_ VPWR VGND sg13g2_xnor2_1
X_4113_ falu_i.falutop.div_inst.b1\[2\] falu_i.falutop.div_inst.acc\[2\] _1115_ VPWR
+ VGND sg13g2_nor2b_1
XFILLER_25_1027 VPWR VGND sg13g2_fill_2
XFILLER_37_531 VPWR VGND sg13g2_fill_2
X_4044_ _1067_ _2441_ _1049_ VPWR VGND sg13g2_nand2b_1
X_4946_ _1840_ _1889_ _0304_ VPWR VGND sg13g2_nor2_1
XFILLER_21_910 VPWR VGND sg13g2_decap_8
X_4877_ _1819_ _1821_ _1822_ VPWR VGND sg13g2_nor2_1
XFILLER_20_420 VPWR VGND sg13g2_fill_2
XFILLER_20_431 VPWR VGND sg13g2_fill_1
X_3828_ VGND VPWR _2211_ net642 _0133_ _0942_ sg13g2_a21oi_1
XFILLER_21_987 VPWR VGND sg13g2_decap_8
XFILLER_4_619 VPWR VGND sg13g2_decap_4
X_3759_ net883 _0906_ _0907_ VPWR VGND sg13g2_and2_1
X_5317__67 VPWR VGND net67 sg13g2_tiehi
X_5332__37 VPWR VGND net37 sg13g2_tiehi
X_5480__325 VPWR VGND net325 sg13g2_tiehi
X_5429_ net176 VGND VPWR _0188_ ppwm_i.u_ppwm.u_mem.memory\[88\] clknet_leaf_32_clk
+ sg13g2_dfrbpq_1
XFILLER_0_869 VPWR VGND sg13g2_decap_8
XFILLER_47_328 VPWR VGND sg13g2_decap_4
XFILLER_28_520 VPWR VGND sg13g2_decap_4
XFILLER_16_737 VPWR VGND sg13g2_decap_8
XFILLER_15_236 VPWR VGND sg13g2_decap_4
X_5339__372 VPWR VGND net372 sg13g2_tiehi
XFILLER_24_781 VPWR VGND sg13g2_decap_8
XFILLER_12_965 VPWR VGND sg13g2_decap_8
XFILLER_23_72 VPWR VGND sg13g2_fill_2
XFILLER_8_958 VPWR VGND sg13g2_decap_8
XFILLER_7_446 VPWR VGND sg13g2_decap_8
XFILLER_48_1005 VPWR VGND sg13g2_decap_8
XFILLER_3_674 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_46_394 VPWR VGND sg13g2_fill_1
XFILLER_46_372 VPWR VGND sg13g2_fill_2
XFILLER_19_597 VPWR VGND sg13g2_decap_8
X_4800_ _1745_ _1742_ _1746_ VPWR VGND sg13g2_xor2_1
X_2992_ VPWR _2346_ _2345_ VGND sg13g2_inv_1
XFILLER_15_770 VPWR VGND sg13g2_decap_8
X_4731_ _1565_ _1638_ _1678_ VPWR VGND _1494_ sg13g2_nand3b_1
XFILLER_9_96 VPWR VGND sg13g2_decap_4
X_4662_ _1272_ _1609_ _1610_ VPWR VGND sg13g2_nor2b_1
X_3613_ net601 VPWR _0781_ VGND ppwm_i.u_ppwm.pwm_value\[7\] ppwm_i.u_ppwm.pwm_value\[6\]
+ sg13g2_o21ai_1
X_4593_ _1475_ VPWR _1542_ VGND _1462_ _1476_ sg13g2_o21ai_1
X_3544_ VGND VPWR _0651_ _0695_ _0716_ net574 sg13g2_a21oi_1
X_3475_ _2251_ net598 _0650_ VPWR VGND sg13g2_nor2_1
XFILLER_9_1021 VPWR VGND sg13g2_decap_8
X_5214_ _2125_ falu_i.falutop.data_in\[6\] _2127_ VPWR VGND sg13g2_xor2_1
X_5282__132 VPWR VGND net132 sg13g2_tiehi
X_5145_ _2066_ _2082_ _2083_ VPWR VGND sg13g2_nor2_1
XFILLER_28_28 VPWR VGND sg13g2_decap_8
X_5076_ VPWR VGND net638 net630 _2016_ net614 _2017_ _2013_ sg13g2_a221oi_1
X_4027_ net459 net1015 _2442_ _1054_ VPWR VGND sg13g2_mux2_1
XFILLER_37_383 VPWR VGND sg13g2_fill_1
XFILLER_37_361 VPWR VGND sg13g2_fill_2
XFILLER_25_512 VPWR VGND sg13g2_decap_4
X_4929_ VGND VPWR _1870_ _1871_ _1873_ _1843_ sg13g2_a21oi_1
XFILLER_0_611 VPWR VGND sg13g2_fill_2
XFILLER_0_633 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_0_699 VPWR VGND sg13g2_decap_8
XFILLER_28_372 VPWR VGND sg13g2_decap_8
X_5487__309 VPWR VGND net309 sg13g2_tiehi
XFILLER_15_1015 VPWR VGND sg13g2_decap_8
XFILLER_8_755 VPWR VGND sg13g2_fill_2
XFILLER_12_784 VPWR VGND sg13g2_fill_1
XFILLER_8_777 VPWR VGND sg13g2_fill_1
XFILLER_4_950 VPWR VGND sg13g2_decap_8
X_3260_ net1129 _0445_ net974 _0449_ VPWR VGND sg13g2_nand3_1
XFILLER_22_4 VPWR VGND sg13g2_decap_8
X_3191_ _0402_ net1118 _0035_ VPWR VGND sg13g2_nor2_1
XFILLER_26_309 VPWR VGND sg13g2_fill_1
XFILLER_34_320 VPWR VGND sg13g2_fill_2
XFILLER_35_843 VPWR VGND sg13g2_fill_1
X_2975_ _2328_ VPWR _2329_ VGND _2316_ _2321_ sg13g2_o21ai_1
X_4714_ _1661_ _1658_ _1659_ VPWR VGND sg13g2_xnor2_1
X_4645_ VGND VPWR net739 net715 _1593_ net750 sg13g2_a21oi_1
X_4576_ VGND VPWR _1524_ _1525_ _1526_ _1406_ sg13g2_a21oi_1
X_3527_ _0699_ VPWR _0700_ VGND _2245_ net597 sg13g2_o21ai_1
X_3458_ _0634_ net611 _0633_ VPWR VGND sg13g2_nand2_1
X_3389_ net782 _2267_ _0563_ _0567_ VPWR VGND sg13g2_nor3_1
X_5128_ VGND VPWR _2053_ _2065_ _2067_ _2066_ sg13g2_a21oi_1
XFILLER_44_106 VPWR VGND sg13g2_decap_8
X_5059_ _2000_ _1991_ _1998_ VPWR VGND sg13g2_xnor2_1
X_5516__221 VPWR VGND net221 sg13g2_tiehi
XFILLER_40_301 VPWR VGND sg13g2_fill_1
XFILLER_40_356 VPWR VGND sg13g2_fill_2
XFILLER_4_202 VPWR VGND sg13g2_decap_8
XFILLER_5_769 VPWR VGND sg13g2_decap_4
XFILLER_20_40 VPWR VGND sg13g2_fill_2
XFILLER_1_931 VPWR VGND sg13g2_decap_8
XFILLER_49_957 VPWR VGND sg13g2_decap_8
Xhold71 ppwm_i.u_ppwm.u_mem.memory\[53\] VPWR VGND net443 sg13g2_dlygate4sd3_1
Xhold60 falu_i.falutop.div_inst.quo\[5\] VPWR VGND net432 sg13g2_dlygate4sd3_1
Xhold82 ppwm_i.u_ppwm.u_mem.memory\[104\] VPWR VGND net454 sg13g2_dlygate4sd3_1
Xhold93 falu_i.falutop.div_inst.a\[5\] VPWR VGND net465 sg13g2_dlygate4sd3_1
XFILLER_44_684 VPWR VGND sg13g2_decap_8
XFILLER_17_876 VPWR VGND sg13g2_decap_8
XFILLER_44_695 VPWR VGND sg13g2_fill_2
XFILLER_43_183 VPWR VGND sg13g2_decap_8
XFILLER_16_386 VPWR VGND sg13g2_decap_4
XFILLER_12_570 VPWR VGND sg13g2_decap_4
XFILLER_8_552 VPWR VGND sg13g2_decap_4
X_4430_ _1382_ _1324_ _1231_ _1322_ _1235_ VPWR VGND sg13g2_a22oi_1
XFILLER_6_53 VPWR VGND sg13g2_fill_1
XFILLER_6_97 VPWR VGND sg13g2_decap_4
X_4361_ _1314_ _1305_ VPWR VGND _1260_ sg13g2_nand2b_2
XFILLER_4_791 VPWR VGND sg13g2_decap_4
X_4292_ net717 net747 _1245_ VPWR VGND sg13g2_nor2_1
X_3312_ net419 net799 _0493_ VPWR VGND sg13g2_nor2_1
X_3243_ VGND VPWR ppwm_i.u_ppwm.global_counter\[7\] _0435_ _0438_ net553 sg13g2_a21oi_1
X_3174_ VGND VPWR _2283_ net682 _0029_ _0392_ sg13g2_a21oi_1
X_5498__279 VPWR VGND net279 sg13g2_tiehi
XFILLER_23_835 VPWR VGND sg13g2_decap_8
XFILLER_22_367 VPWR VGND sg13g2_fill_2
X_2958_ net792 net794 _2312_ VPWR VGND sg13g2_nor2b_2
X_2889_ _2243_ ppwm_i.u_ppwm.pwm_value\[9\] VPWR VGND sg13g2_inv_2
X_4628_ VPWR VGND _1239_ _1574_ _1383_ _1236_ _1577_ _1319_ sg13g2_a221oi_1
Xhold530 _0076_ VPWR VGND net1182 sg13g2_dlygate4sd3_1
Xhold541 ppwm_i.u_ppwm.pc\[2\] VPWR VGND net1193 sg13g2_dlygate4sd3_1
X_4559_ _1314_ VPWR _1509_ VGND net734 net759 sg13g2_o21ai_1
XFILLER_46_916 VPWR VGND sg13g2_decap_8
XFILLER_17_117 VPWR VGND sg13g2_fill_1
XFILLER_26_640 VPWR VGND sg13g2_fill_2
X_5373__306 VPWR VGND net306 sg13g2_tiehi
XFILLER_14_802 VPWR VGND sg13g2_fill_2
XFILLER_14_824 VPWR VGND sg13g2_decap_8
XFILLER_25_150 VPWR VGND sg13g2_fill_2
XFILLER_26_662 VPWR VGND sg13g2_decap_8
XFILLER_41_632 VPWR VGND sg13g2_fill_2
XFILLER_13_323 VPWR VGND sg13g2_fill_2
XFILLER_41_698 VPWR VGND sg13g2_fill_1
XFILLER_12_1007 VPWR VGND sg13g2_decap_8
XFILLER_5_533 VPWR VGND sg13g2_fill_1
XFILLER_31_94 VPWR VGND sg13g2_fill_1
X_5419__214 VPWR VGND net214 sg13g2_tiehi
XFILLER_45_971 VPWR VGND sg13g2_decap_8
X_3930_ VGND VPWR _2174_ net673 _0184_ _0993_ sg13g2_a21oi_1
XFILLER_17_695 VPWR VGND sg13g2_decap_4
X_3861_ net831 VPWR _0959_ VGND ppwm_i.u_ppwm.u_mem.memory\[51\] net643 sg13g2_o21ai_1
XFILLER_32_643 VPWR VGND sg13g2_fill_2
X_3792_ VGND VPWR _2224_ net644 _0115_ _0924_ sg13g2_a21oi_1
X_2812_ VPWR _2166_ net562 VGND sg13g2_inv_1
X_5531_ net137 VGND VPWR net857 falu_i.falutop.div_inst.acc\[4\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_8_382 VPWR VGND sg13g2_fill_2
X_5430__171 VPWR VGND net171 sg13g2_tiehi
X_5462_ net38 VGND VPWR _0221_ falu_i.falutop.i2c_inst.state\[1\] clknet_leaf_9_clk
+ sg13g2_dfrbpq_2
X_5393_ net266 VGND VPWR net444 ppwm_i.u_ppwm.u_mem.memory\[52\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4413_ _1365_ _1364_ _1299_ VPWR VGND sg13g2_nand2b_1
X_4344_ _1296_ VPWR _1297_ VGND net707 net587 sg13g2_o21ai_1
X_4275_ _1228_ net736 net765 VPWR VGND sg13g2_nand2_2
XFILLER_39_231 VPWR VGND sg13g2_fill_1
X_3226_ VGND VPWR _0427_ _0425_ _2272_ sg13g2_or2_1
XFILLER_39_286 VPWR VGND sg13g2_fill_1
X_3157_ net820 VPWR _0383_ VGND net1044 _0382_ sg13g2_o21ai_1
XFILLER_28_938 VPWR VGND sg13g2_decap_8
XFILLER_43_919 VPWR VGND sg13g2_decap_8
X_3088_ falu_i.falutop.i2c_inst.counter\[1\] net1045 _2438_ VPWR VGND sg13g2_nor2_2
XFILLER_22_120 VPWR VGND sg13g2_fill_1
XFILLER_23_665 VPWR VGND sg13g2_fill_2
XFILLER_7_809 VPWR VGND sg13g2_fill_1
XFILLER_2_514 VPWR VGND sg13g2_decap_8
Xhold371 _0295_ VPWR VGND net1023 sg13g2_dlygate4sd3_1
Xhold360 _0216_ VPWR VGND net1012 sg13g2_dlygate4sd3_1
Xhold382 _0303_ VPWR VGND net1034 sg13g2_dlygate4sd3_1
Xhold393 falu_i.falutop.i2c_inst.counter\[0\] VPWR VGND net1045 sg13g2_dlygate4sd3_1
Xfanout840 net841 net840 VPWR VGND sg13g2_buf_8
XFILLER_19_905 VPWR VGND sg13g2_decap_8
XFILLER_45_267 VPWR VGND sg13g2_fill_2
XFILLER_45_256 VPWR VGND sg13g2_fill_2
XFILLER_14_632 VPWR VGND sg13g2_decap_8
XFILLER_42_952 VPWR VGND sg13g2_decap_8
XFILLER_6_864 VPWR VGND sg13g2_decap_8
X_4060_ net901 falu_i.falutop.data_in\[1\] net684 _0229_ VPWR VGND sg13g2_mux2_1
XFILLER_49_584 VPWR VGND sg13g2_decap_4
X_3011_ net691 ppwm_i.u_ppwm.u_mem.memory\[69\] net789 _2365_ VPWR VGND sg13g2_a21o_1
XFILLER_37_702 VPWR VGND sg13g2_decap_4
X_4962_ VGND VPWR net718 _1803_ _1905_ _1904_ sg13g2_a21oi_1
X_3913_ net839 VPWR _0985_ VGND net404 net676 sg13g2_o21ai_1
X_4893_ VPWR VGND _1837_ net630 net614 falu_i.falutop.div_inst.rem\[0\] _1838_ net638
+ sg13g2_a221oi_1
XFILLER_33_974 VPWR VGND sg13g2_decap_8
X_3844_ VGND VPWR _2206_ net656 _0141_ _0950_ sg13g2_a21oi_1
XFILLER_20_635 VPWR VGND sg13g2_decap_4
X_5329__43 VPWR VGND net43 sg13g2_tiehi
XFILLER_20_668 VPWR VGND sg13g2_decap_8
X_3775_ net835 VPWR _0916_ VGND net451 net662 sg13g2_o21ai_1
X_5514_ net229 VGND VPWR net1099 falu_i.falutop.div_inst.rem\[1\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_5445_ net110 VGND VPWR _0204_ ppwm_i.u_ppwm.u_mem.memory\[104\] clknet_leaf_30_clk
+ sg13g2_dfrbpq_2
X_5376_ net300 VGND VPWR net473 ppwm_i.u_ppwm.u_mem.memory\[35\] clknet_leaf_22_clk
+ sg13g2_dfrbpq_1
X_4327_ net772 _1279_ _1280_ VPWR VGND sg13g2_nor2_1
XFILLER_41_1011 VPWR VGND sg13g2_decap_8
X_4258_ _1212_ VPWR _0293_ VGND _1098_ _1179_ sg13g2_o21ai_1
X_3209_ VGND VPWR _0416_ _0415_ net1177 sg13g2_or2_1
X_4189_ _1162_ VPWR _1163_ VGND net489 _1132_ sg13g2_o21ai_1
XFILLER_24_963 VPWR VGND sg13g2_decap_8
XFILLER_10_134 VPWR VGND sg13g2_fill_2
XFILLER_11_657 VPWR VGND sg13g2_decap_8
XFILLER_23_495 VPWR VGND sg13g2_decap_8
XFILLER_3_889 VPWR VGND sg13g2_decap_8
XFILLER_2_355 VPWR VGND sg13g2_fill_1
Xhold190 ppwm_i.u_ppwm.u_mem.memory\[98\] VPWR VGND net562 sg13g2_dlygate4sd3_1
Xfanout670 net671 net670 VPWR VGND sg13g2_buf_8
Xfanout681 net683 net681 VPWR VGND sg13g2_buf_8
Xfanout692 _2311_ net692 VPWR VGND sg13g2_buf_8
XFILLER_37_71 VPWR VGND sg13g2_fill_2
XFILLER_33_215 VPWR VGND sg13g2_fill_1
XFILLER_15_952 VPWR VGND sg13g2_decap_8
XFILLER_42_793 VPWR VGND sg13g2_decap_8
XFILLER_41_281 VPWR VGND sg13g2_fill_2
XFILLER_30_944 VPWR VGND sg13g2_decap_8
X_3560_ _0729_ VPWR _0731_ VGND _0708_ _0712_ sg13g2_o21ai_1
X_5269__158 VPWR VGND net158 sg13g2_tiehi
XFILLER_6_683 VPWR VGND sg13g2_decap_4
X_5230_ _2091_ net776 _2138_ VPWR VGND sg13g2_nor2b_1
X_3491_ net573 _0660_ _0664_ _0665_ _0666_ VPWR VGND sg13g2_nor4_1
X_5161_ falu_i.falutop.data_in\[3\] _2096_ _2097_ VPWR VGND sg13g2_nor2b_1
X_5092_ _2032_ _1994_ _2031_ VPWR VGND sg13g2_xnor2_1
X_4112_ falu_i.falutop.div_inst.b1\[3\] falu_i.falutop.div_inst.acc\[3\] _1114_ VPWR
+ VGND sg13g2_nor2b_1
X_4043_ net797 _1066_ _0224_ VPWR VGND sg13g2_nor2_1
XFILLER_49_392 VPWR VGND sg13g2_decap_4
XFILLER_24_215 VPWR VGND sg13g2_decap_4
XFILLER_25_749 VPWR VGND sg13g2_decap_8
X_4945_ VPWR VGND _1888_ net630 _1886_ net614 _1889_ _1885_ sg13g2_a221oi_1
X_4876_ VGND VPWR _1817_ _1818_ _1821_ _1800_ sg13g2_a21oi_1
XFILLER_20_410 VPWR VGND sg13g2_fill_1
XFILLER_21_966 VPWR VGND sg13g2_decap_8
XFILLER_32_281 VPWR VGND sg13g2_decap_4
X_3827_ net826 VPWR _0942_ VGND ppwm_i.u_ppwm.u_mem.memory\[34\] net642 sg13g2_o21ai_1
XFILLER_20_498 VPWR VGND sg13g2_decap_4
X_3758_ ppwm_i.u_ppwm.u_mem.clk_prog_sync3 net375 _0906_ VPWR VGND sg13g2_nor2b_2
X_3689_ _0618_ _0850_ _0851_ VPWR VGND sg13g2_nor2_1
X_5428_ net180 VGND VPWR net519 ppwm_i.u_ppwm.u_mem.memory\[87\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_0_848 VPWR VGND sg13g2_decap_8
X_5359_ net334 VGND VPWR _0118_ ppwm_i.u_ppwm.u_mem.memory\[18\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
XFILLER_28_576 VPWR VGND sg13g2_fill_2
XFILLER_24_760 VPWR VGND sg13g2_decap_8
XFILLER_12_944 VPWR VGND sg13g2_decap_8
XFILLER_8_937 VPWR VGND sg13g2_decap_8
XFILLER_11_498 VPWR VGND sg13g2_decap_8
XFILLER_48_1028 VPWR VGND sg13g2_fill_1
XFILLER_0_77 VPWR VGND sg13g2_decap_8
X_2991_ _2329_ _2344_ _2345_ VPWR VGND sg13g2_and2_1
X_4730_ VPWR VGND net631 _1676_ _1668_ net616 _1677_ _1666_ sg13g2_a221oi_1
XFILLER_9_64 VPWR VGND sg13g2_fill_1
X_4661_ _1270_ _1271_ _1217_ _1609_ VPWR VGND sg13g2_nand3_1
X_3612_ _0729_ _0746_ _0712_ _0780_ VPWR VGND _0765_ sg13g2_nand4_1
XFILLER_31_1010 VPWR VGND sg13g2_decap_8
X_4592_ _1541_ _1527_ _1539_ VPWR VGND sg13g2_xnor2_1
X_3543_ _0635_ _0714_ _0715_ VPWR VGND sg13g2_nor2_1
XFILLER_43_0 VPWR VGND sg13g2_decap_4
X_3474_ VGND VPWR _0649_ _0620_ _2419_ sg13g2_or2_1
XFILLER_9_1000 VPWR VGND sg13g2_decap_8
X_5213_ net920 net623 _2126_ VPWR VGND sg13g2_nor2_1
X_5144_ _2081_ VPWR _2082_ VGND _2063_ _2064_ sg13g2_o21ai_1
XFILLER_29_318 VPWR VGND sg13g2_decap_8
X_5075_ _2014_ _2015_ _2016_ VPWR VGND sg13g2_and2_1
X_4026_ _1051_ VPWR _1053_ VGND _1049_ _1052_ sg13g2_o21ai_1
XFILLER_38_885 VPWR VGND sg13g2_fill_1
X_4928_ _1870_ _1871_ _1843_ _1872_ VPWR VGND sg13g2_nand3_1
X_4859_ net768 net752 net711 _1804_ VPWR VGND sg13g2_nand3_1
Xclkbuf_3_0__f_clk clknet_0_clk clknet_3_0__leaf_clk VPWR VGND sg13g2_buf_8
XFILLER_48_627 VPWR VGND sg13g2_fill_1
XFILLER_28_351 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_16_535 VPWR VGND sg13g2_fill_1
XFILLER_16_546 VPWR VGND sg13g2_decap_8
XFILLER_43_387 VPWR VGND sg13g2_fill_2
XFILLER_8_701 VPWR VGND sg13g2_fill_2
XFILLER_34_94 VPWR VGND sg13g2_fill_1
XFILLER_3_494 VPWR VGND sg13g2_fill_2
X_3190_ net808 VPWR _0403_ VGND net1117 _0400_ sg13g2_o21ai_1
XFILLER_15_4 VPWR VGND sg13g2_fill_1
XFILLER_19_351 VPWR VGND sg13g2_fill_2
XFILLER_34_365 VPWR VGND sg13g2_fill_2
XFILLER_34_376 VPWR VGND sg13g2_decap_4
X_2974_ _2327_ VPWR _2328_ VGND _2324_ _2326_ sg13g2_o21ai_1
X_4713_ _1658_ _1659_ _1660_ VPWR VGND sg13g2_nor2_1
X_4644_ _1592_ net739 net715 net750 VPWR VGND sg13g2_and3_1
X_4575_ _1525_ _1523_ net947 VPWR VGND sg13g2_nand2b_1
X_3526_ _0699_ ppwm_i.u_ppwm.u_ex.reg_value_q\[7\] net596 VPWR VGND sg13g2_nand2_1
X_3457_ VGND VPWR _0632_ _0633_ net595 _2241_ sg13g2_a21oi_2
X_3388_ _0566_ _2235_ ppwm_i.u_ppwm.global_counter\[9\] VPWR VGND sg13g2_nand2_1
X_5127_ net615 VPWR _2066_ VGND _2053_ _2065_ sg13g2_o21ai_1
X_5058_ _1991_ _1998_ _1999_ VPWR VGND sg13g2_nor2_1
X_4009_ VGND VPWR _1022_ _1039_ _1040_ net796 sg13g2_a21oi_1
XFILLER_38_1027 VPWR VGND sg13g2_fill_2
XFILLER_38_1016 VPWR VGND sg13g2_decap_8
XFILLER_13_505 VPWR VGND sg13g2_fill_1
XFILLER_13_516 VPWR VGND sg13g2_decap_4
XFILLER_26_888 VPWR VGND sg13g2_decap_8
XFILLER_40_379 VPWR VGND sg13g2_decap_8
XFILLER_21_582 VPWR VGND sg13g2_fill_1
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_0_453 VPWR VGND sg13g2_decap_4
XFILLER_1_987 VPWR VGND sg13g2_decap_8
XFILLER_49_936 VPWR VGND sg13g2_decap_8
Xhold50 ppwm_i.u_ppwm.u_mem.memory\[39\] VPWR VGND net422 sg13g2_dlygate4sd3_1
XFILLER_0_497 VPWR VGND sg13g2_decap_8
Xhold72 _0152_ VPWR VGND net444 sg13g2_dlygate4sd3_1
Xhold83 ppwm_i.u_ppwm.u_mem.memory\[40\] VPWR VGND net455 sg13g2_dlygate4sd3_1
Xhold61 _0284_ VPWR VGND net433 sg13g2_dlygate4sd3_1
Xhold94 _0341_ VPWR VGND net466 sg13g2_dlygate4sd3_1
XFILLER_29_660 VPWR VGND sg13g2_fill_1
XFILLER_29_671 VPWR VGND sg13g2_decap_8
XFILLER_17_855 VPWR VGND sg13g2_decap_8
XFILLER_43_151 VPWR VGND sg13g2_fill_2
XFILLER_6_10 VPWR VGND sg13g2_decap_8
X_4360_ _1260_ _1305_ _1313_ VPWR VGND sg13g2_nor2b_1
X_3311_ _0491_ VPWR _0492_ VGND _0479_ _0488_ sg13g2_o21ai_1
X_4291_ _1244_ net720 net747 VPWR VGND sg13g2_nand2_2
X_3242_ net796 net1093 _0052_ VPWR VGND sg13g2_nor2_1
X_3173_ net810 VPWR _0392_ VGND ppwm_i.u_ppwm.pwm_value\[5\] net682 sg13g2_o21ai_1
XFILLER_6_1025 VPWR VGND sg13g2_decap_4
XFILLER_48_991 VPWR VGND sg13g2_decap_8
XFILLER_23_814 VPWR VGND sg13g2_decap_8
XFILLER_22_302 VPWR VGND sg13g2_decap_4
XFILLER_41_18 VPWR VGND sg13g2_fill_2
X_2957_ net794 net792 _2311_ VPWR VGND sg13g2_nor2b_2
X_2888_ net1144 _2242_ VPWR VGND sg13g2_inv_4
X_4627_ _1575_ VPWR _1576_ VGND _1239_ _1323_ sg13g2_o21ai_1
Xhold520 ppwm_i.u_ppwm.u_ex.reg_value_q\[6\] VPWR VGND net1172 sg13g2_dlygate4sd3_1
Xhold542 ppwm_i.u_ppwm.u_ex.reg_value_q\[8\] VPWR VGND net1194 sg13g2_dlygate4sd3_1
Xhold531 ppwm_i.u_ppwm.u_ex.reg_value_q\[4\] VPWR VGND net1183 sg13g2_dlygate4sd3_1
X_4558_ _1506_ _1225_ _1508_ VPWR VGND sg13g2_xor2_1
X_4489_ _1440_ _1229_ _1267_ VPWR VGND sg13g2_nand2_1
X_3509_ net577 VPWR _0683_ VGND ppwm_i.u_ppwm.u_ex.reg_value_q\[2\] net588 sg13g2_o21ai_1
XFILLER_39_980 VPWR VGND sg13g2_decap_8
XFILLER_18_619 VPWR VGND sg13g2_fill_1
XFILLER_45_449 VPWR VGND sg13g2_fill_2
Xclkbuf_leaf_37_clk clknet_3_5__leaf_clk clknet_leaf_37_clk VPWR VGND sg13g2_buf_8
XFILLER_26_652 VPWR VGND sg13g2_fill_1
XFILLER_13_313 VPWR VGND sg13g2_fill_1
XFILLER_25_184 VPWR VGND sg13g2_fill_1
XFILLER_13_335 VPWR VGND sg13g2_decap_8
XFILLER_13_346 VPWR VGND sg13g2_fill_1
XFILLER_22_880 VPWR VGND sg13g2_decap_8
X_5447__102 VPWR VGND net102 sg13g2_tiehi
XFILLER_31_73 VPWR VGND sg13g2_fill_2
XFILLER_1_751 VPWR VGND sg13g2_decap_4
XFILLER_49_711 VPWR VGND sg13g2_decap_8
XFILLER_0_261 VPWR VGND sg13g2_fill_2
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_49_777 VPWR VGND sg13g2_decap_8
XFILLER_49_788 VPWR VGND sg13g2_fill_2
XFILLER_36_405 VPWR VGND sg13g2_decap_4
XFILLER_45_950 VPWR VGND sg13g2_decap_8
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk clknet_leaf_28_clk VPWR VGND sg13g2_buf_8
XFILLER_44_471 VPWR VGND sg13g2_fill_2
X_3860_ VGND VPWR _2200_ net664 _0149_ _0958_ sg13g2_a21oi_1
XFILLER_13_880 VPWR VGND sg13g2_decap_8
XFILLER_20_839 VPWR VGND sg13g2_decap_8
X_3791_ net828 VPWR _0924_ VGND net515 net644 sg13g2_o21ai_1
X_2811_ VPWR _2165_ net537 VGND sg13g2_inv_1
X_5530_ net145 VGND VPWR net495 falu_i.falutop.div_inst.acc\[3\] clknet_leaf_0_clk
+ sg13g2_dfrbpq_2
XFILLER_9_895 VPWR VGND sg13g2_decap_8
X_5461_ net42 VGND VPWR net460 falu_i.falutop.i2c_inst.state\[0\] clknet_leaf_10_clk
+ sg13g2_dfrbpq_2
X_4412_ _1363_ net743 _1364_ VPWR VGND net587 sg13g2_nand3b_1
X_5392_ net268 VGND VPWR net916 ppwm_i.u_ppwm.u_mem.memory\[51\] clknet_leaf_25_clk
+ sg13g2_dfrbpq_1
X_4343_ _1296_ net743 net587 VPWR VGND sg13g2_nand2_1
XFILLER_28_1015 VPWR VGND sg13g2_decap_8
X_4274_ net737 net763 _1227_ VPWR VGND sg13g2_and2_1
X_3225_ net943 _0426_ _0046_ VPWR VGND sg13g2_nor2_1
X_3156_ _2431_ _0344_ _0382_ VPWR VGND sg13g2_nor2_1
XFILLER_28_917 VPWR VGND sg13g2_decap_8
XFILLER_36_18 VPWR VGND sg13g2_fill_2
XFILLER_43_909 VPWR VGND sg13g2_fill_1
X_5279__138 VPWR VGND net138 sg13g2_tiehi
X_3087_ _2437_ _2430_ VPWR VGND net1150 sg13g2_nand2b_2
Xclkbuf_leaf_19_clk clknet_3_4__leaf_clk clknet_leaf_19_clk VPWR VGND sg13g2_buf_8
XFILLER_36_983 VPWR VGND sg13g2_decap_8
XFILLER_11_806 VPWR VGND sg13g2_decap_4
XFILLER_23_644 VPWR VGND sg13g2_decap_8
XFILLER_35_1019 VPWR VGND sg13g2_decap_8
XFILLER_11_839 VPWR VGND sg13g2_decap_8
XFILLER_22_154 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_fill_1
XFILLER_23_677 VPWR VGND sg13g2_fill_2
X_3989_ net652 _1021_ net1152 _1024_ VPWR VGND sg13g2_nand3_1
XFILLER_2_537 VPWR VGND sg13g2_fill_1
Xhold361 falu_i.falutop.i2c_inst.counter\[2\] VPWR VGND net1013 sg13g2_dlygate4sd3_1
Xhold350 _2447_ VPWR VGND net1002 sg13g2_dlygate4sd3_1
Xhold372 ppwm_i.u_ppwm.u_pwm.counter\[9\] VPWR VGND net1024 sg13g2_dlygate4sd3_1
Xhold383 falu_i.falutop.i2c_inst.result\[13\] VPWR VGND net1035 sg13g2_dlygate4sd3_1
Xhold394 _0343_ VPWR VGND net1046 sg13g2_dlygate4sd3_1
Xfanout841 net842 net841 VPWR VGND sg13g2_buf_8
Xfanout830 net831 net830 VPWR VGND sg13g2_buf_8
XFILLER_26_51 VPWR VGND sg13g2_fill_1
XFILLER_42_931 VPWR VGND sg13g2_decap_8
XFILLER_27_994 VPWR VGND sg13g2_decap_8
XFILLER_13_132 VPWR VGND sg13g2_decap_8
XFILLER_14_666 VPWR VGND sg13g2_decap_8
XFILLER_9_114 VPWR VGND sg13g2_fill_1
XFILLER_14_677 VPWR VGND sg13g2_fill_2
XFILLER_6_810 VPWR VGND sg13g2_decap_4
XFILLER_6_843 VPWR VGND sg13g2_decap_8
XFILLER_10_894 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_3_99 VPWR VGND sg13g2_decap_8
X_3010_ _2364_ ppwm_i.u_ppwm.u_mem.memory\[83\] net702 VPWR VGND sg13g2_nand2_1
XFILLER_37_758 VPWR VGND sg13g2_decap_8
X_4961_ _1904_ net753 net718 net768 net711 VPWR VGND sg13g2_a22oi_1
X_3912_ VGND VPWR _2182_ net649 _0175_ _0984_ sg13g2_a21oi_1
X_4892_ _1831_ _1834_ _1787_ _1837_ VPWR VGND _1836_ sg13g2_nand4_1
XFILLER_33_953 VPWR VGND sg13g2_decap_8
X_3843_ net825 VPWR _0950_ VGND ppwm_i.u_ppwm.u_mem.memory\[41\] net656 sg13g2_o21ai_1
X_3774_ VGND VPWR _2230_ net654 _0106_ _0915_ sg13g2_a21oi_1
X_5513_ net233 VGND VPWR _0272_ falu_i.falutop.div_inst.rem\[0\] clknet_leaf_1_clk
+ sg13g2_dfrbpq_2
X_5444_ net114 VGND VPWR _0203_ ppwm_i.u_ppwm.u_mem.memory\[103\] clknet_leaf_31_clk
+ sg13g2_dfrbpq_1
Xclkbuf_leaf_8_clk clknet_3_2__leaf_clk clknet_leaf_8_clk VPWR VGND sg13g2_buf_8
X_5375_ net302 VGND VPWR _0134_ ppwm_i.u_ppwm.u_mem.memory\[34\] clknet_leaf_23_clk
+ sg13g2_dfrbpq_1
X_4326_ _1279_ falu_i.falutop.alu_inst.op\[1\] _2298_ VPWR VGND sg13g2_nand2_2
X_4257_ _1212_ net485 net607 VPWR VGND sg13g2_nand2_1
X_3208_ net796 net1067 _0415_ _0040_ VPWR VGND sg13g2_nor3_1
X_4188_ _1162_ net568 _1161_ VPWR VGND sg13g2_nand2_1
X_3139_ net816 VPWR _0371_ VGND net926 _0370_ sg13g2_o21ai_1
XFILLER_27_202 VPWR VGND sg13g2_fill_1
XFILLER_16_909 VPWR VGND sg13g2_decap_8
X_5292__113 VPWR VGND net113 sg13g2_tiehi
XFILLER_42_216 VPWR VGND sg13g2_fill_2
XFILLER_42_249 VPWR VGND sg13g2_decap_8
XFILLER_24_942 VPWR VGND sg13g2_decap_8
XFILLER_11_603 VPWR VGND sg13g2_fill_2
XFILLER_11_636 VPWR VGND sg13g2_fill_2
XFILLER_11_647 VPWR VGND sg13g2_decap_4
XFILLER_7_629 VPWR VGND sg13g2_fill_1
Xhold180 _0177_ VPWR VGND net552 sg13g2_dlygate4sd3_1
XFILLER_3_868 VPWR VGND sg13g2_decap_8
Xhold191 ppwm_i.u_ppwm.u_mem.memory\[77\] VPWR VGND net843 sg13g2_dlygate4sd3_1
Xfanout660 net663 net660 VPWR VGND sg13g2_buf_1
X_5305__223 VPWR VGND net223 sg13g2_tiehi
Xfanout682 net683 net682 VPWR VGND sg13g2_buf_8
Xfanout671 net679 net671 VPWR VGND sg13g2_buf_8
Xfanout693 _2311_ net693 VPWR VGND sg13g2_buf_2
XFILLER_46_544 VPWR VGND sg13g2_decap_8
XFILLER_37_61 VPWR VGND sg13g2_fill_2
XFILLER_34_706 VPWR VGND sg13g2_fill_2
XFILLER_46_588 VPWR VGND sg13g2_fill_2
XFILLER_15_931 VPWR VGND sg13g2_decap_8
XFILLER_42_761 VPWR VGND sg13g2_decap_4
XFILLER_30_923 VPWR VGND sg13g2_decap_8
XFILLER_41_293 VPWR VGND sg13g2_decap_8
X_3490_ _2381_ _2388_ _0637_ _0665_ VPWR VGND sg13g2_nor3_1
X_5160_ falu_i.falutop.data_in\[0\] falu_i.falutop.data_in\[1\] falu_i.falutop.data_in\[2\]
+ _2096_ VPWR VGND sg13g2_nor3_1
X_5091_ _2031_ _2025_ _2029_ VPWR VGND sg13g2_xnor2_1
XFILLER_2_890 VPWR VGND sg13g2_decap_8
X_4111_ falu_i.falutop.div_inst.b1\[4\] falu_i.falutop.div_inst.acc\[4\] _1113_ VPWR
+ VGND sg13g2_nor2b_1
X_4042_ _1065_ VPWR _1066_ VGND net1006 _1059_ sg13g2_o21ai_1
XFILLER_37_588 VPWR VGND sg13g2_fill_1
XFILLER_25_728 VPWR VGND sg13g2_decap_8
X_4944_ _1074_ _1887_ _1888_ VPWR VGND sg13g2_nor2_1
XFILLER_24_238 VPWR VGND sg13g2_decap_4
X_4875_ _1817_ _1818_ _1800_ _1820_ VPWR VGND sg13g2_nand3_1
XFILLER_20_422 VPWR VGND sg13g2_fill_1
XFILLER_21_945 VPWR VGND sg13g2_decap_8
X_3826_ VGND VPWR _2211_ net658 _0132_ _0941_ sg13g2_a21oi_1
X_3757_ net807 net4 _0099_ VPWR VGND sg13g2_and2_1
X_3688_ _0848_ _0849_ _0850_ VPWR VGND sg13g2_and2_1
X_5427_ net184 VGND VPWR _0186_ ppwm_i.u_ppwm.u_mem.memory\[86\] clknet_leaf_29_clk
+ sg13g2_dfrbpq_1
XFILLER_0_827 VPWR VGND sg13g2_decap_8
X_5358_ net336 VGND VPWR _0117_ ppwm_i.u_ppwm.u_mem.memory\[17\] clknet_leaf_34_clk
+ sg13g2_dfrbpq_1
X_4309_ _1258_ _1261_ _1257_ _1262_ VPWR VGND sg13g2_nand3_1
X_5289_ net119 VGND VPWR _0051_ ppwm_i.u_ppwm.global_counter\[6\] clknet_leaf_16_clk
+ sg13g2_dfrbpq_1
XFILLER_28_533 VPWR VGND sg13g2_decap_8
XFILLER_28_544 VPWR VGND sg13g2_fill_2
XFILLER_43_547 VPWR VGND sg13g2_fill_1
XFILLER_15_249 VPWR VGND sg13g2_fill_2
XFILLER_12_923 VPWR VGND sg13g2_decap_8
XFILLER_8_916 VPWR VGND sg13g2_decap_8
XFILLER_3_632 VPWR VGND sg13g2_decap_8
XFILLER_47_875 VPWR VGND sg13g2_decap_4
XFILLER_0_1009 VPWR VGND sg13g2_decap_8
XFILLER_47_897 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_19_577 VPWR VGND sg13g2_fill_1
XFILLER_34_525 VPWR VGND sg13g2_decap_4
X_2990_ _2337_ _2334_ _2343_ _2344_ VPWR VGND sg13g2_a21o_2
X_4660_ VGND VPWR _2296_ net565 _1608_ _1607_ sg13g2_a21oi_1
X_3611_ VPWR VGND _0779_ net798 _0769_ _2245_ _0079_ net573 sg13g2_a221oi_1
X_4591_ _1527_ _1539_ _1540_ VPWR VGND sg13g2_nor2b_1
X_3542_ _0714_ net584 _0694_ VPWR VGND sg13g2_nand2_2
XFILLER_7_993 VPWR VGND sg13g2_decap_8
X_3473_ _0624_ _0647_ net609 _0648_ VPWR VGND sg13g2_mux2_1
X_5212_ _2125_ net777 _2099_ VPWR VGND sg13g2_nand2_1
X_5143_ _2081_ _2076_ _2080_ VPWR VGND sg13g2_xnor2_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_5074_ falu_i.falutop.div_inst.rem\[4\] _1973_ net773 _2015_ VPWR VGND sg13g2_nand3_1
XFILLER_37_330 VPWR VGND sg13g2_decap_4
X_4025_ _1052_ net1013 _2438_ VPWR VGND sg13g2_xnor2_1
XFILLER_40_506 VPWR VGND sg13g2_fill_1
X_4927_ _1851_ VPWR _1871_ VGND _1867_ _1869_ sg13g2_o21ai_1
X_4858_ _1803_ net711 net768 net752 VPWR VGND sg13g2_and3_2
X_3809_ net827 VPWR _0933_ VGND net402 net659 sg13g2_o21ai_1
X_4789_ net632 _1383_ _1735_ VPWR VGND sg13g2_nor2_1
XFILLER_28_330 VPWR VGND sg13g2_decap_4
XFILLER_43_333 VPWR VGND sg13g2_fill_2
XFILLER_12_720 VPWR VGND sg13g2_decap_8
XFILLER_11_274 VPWR VGND sg13g2_fill_2
XFILLER_8_757 VPWR VGND sg13g2_fill_1
XFILLER_7_245 VPWR VGND sg13g2_fill_1
XFILLER_4_985 VPWR VGND sg13g2_decap_8
XFILLER_38_116 VPWR VGND sg13g2_fill_1
XFILLER_19_363 VPWR VGND sg13g2_fill_1
XFILLER_35_823 VPWR VGND sg13g2_decap_4
XFILLER_46_193 VPWR VGND sg13g2_fill_2
XFILLER_46_171 VPWR VGND sg13g2_fill_2
XFILLER_22_506 VPWR VGND sg13g2_fill_2
X_2973_ VGND VPWR _2322_ _2323_ _2327_ net787 sg13g2_a21oi_1
XFILLER_22_528 VPWR VGND sg13g2_decap_8
X_4712_ VGND VPWR _1591_ _1599_ _1659_ _1598_ sg13g2_a21oi_1
XFILLER_30_572 VPWR VGND sg13g2_decap_8
XFILLER_30_583 VPWR VGND sg13g2_fill_1
X_4643_ net731 net716 _1591_ VPWR VGND sg13g2_and2_1
X_4574_ _1524_ net947 _1523_ VPWR VGND sg13g2_nand2b_1
X_3525_ net574 _0695_ _0697_ _0698_ VPWR VGND sg13g2_nor3_1
X_3456_ ppwm_i.u_ppwm.pwm_value\[2\] net595 _0632_ VPWR VGND sg13g2_nor2_1
X_3387_ _0562_ _0563_ _0564_ _0565_ VPWR VGND sg13g2_nor3_1
X_5440__130 VPWR VGND net130 sg13g2_tiehi
X_5126_ _2065_ _2063_ _2064_ VPWR VGND sg13g2_xnor2_1
XFILLER_29_116 VPWR VGND sg13g2_fill_1
X_5057_ _1998_ _1939_ _1997_ VPWR VGND sg13g2_xnor2_1
XFILLER_26_823 VPWR VGND sg13g2_fill_2
X_4008_ net883 VPWR _1039_ VGND _1029_ _1038_ sg13g2_o21ai_1
XFILLER_25_344 VPWR VGND sg13g2_fill_1
XFILLER_25_366 VPWR VGND sg13g2_fill_2
XFILLER_26_867 VPWR VGND sg13g2_decap_8
XFILLER_41_837 VPWR VGND sg13g2_fill_1
XFILLER_40_358 VPWR VGND sg13g2_fill_1
X_5486__311 VPWR VGND net311 sg13g2_tiehi
XFILLER_21_594 VPWR VGND sg13g2_decap_4
XFILLER_5_727 VPWR VGND sg13g2_decap_4
XFILLER_20_42 VPWR VGND sg13g2_fill_1
XFILLER_49_915 VPWR VGND sg13g2_decap_8
XFILLER_0_432 VPWR VGND sg13g2_decap_8
XFILLER_1_966 VPWR VGND sg13g2_decap_8
Xhold40 _0281_ VPWR VGND net412 sg13g2_dlygate4sd3_1
XFILLER_0_476 VPWR VGND sg13g2_decap_8
Xhold62 ppwm_i.u_ppwm.u_mem.memory\[49\] VPWR VGND net434 sg13g2_dlygate4sd3_1
Xhold51 _0138_ VPWR VGND net423 sg13g2_dlygate4sd3_1
XFILLER_29_73 VPWR VGND sg13g2_fill_2
Xhold73 ppwm_i.u_ppwm.u_mem.memory\[107\] VPWR VGND net445 sg13g2_dlygate4sd3_1
Xhold84 _0140_ VPWR VGND net456 sg13g2_dlygate4sd3_1
Xhold95 falu_i.falutop.i2c_inst.op\[2\] VPWR VGND net467 sg13g2_dlygate4sd3_1
XFILLER_17_834 VPWR VGND sg13g2_decap_8
X_5462__38 VPWR VGND net38 sg13g2_tiehi
XFILLER_43_130 VPWR VGND sg13g2_fill_2
XFILLER_16_366 VPWR VGND sg13g2_fill_1
XFILLER_32_826 VPWR VGND sg13g2_fill_2
X_3310_ VGND VPWR _0482_ _0487_ _0491_ _0490_ sg13g2_a21oi_1
X_4290_ net717 net747 _1243_ VPWR VGND sg13g2_and2_1
X_3241_ _0437_ net1092 _0435_ VPWR VGND sg13g2_xnor2_1
X_3172_ VGND VPWR _2284_ net681 _0028_ _0391_ sg13g2_a21oi_1
XFILLER_6_1004 VPWR VGND sg13g2_decap_8
XFILLER_48_970 VPWR VGND sg13g2_decap_8
XFILLER_35_631 VPWR VGND sg13g2_fill_2
X_2956_ VGND VPWR _2310_ net794 net792 sg13g2_or2_1
XFILLER_30_391 VPWR VGND sg13g2_decap_8
X_2887_ net1143 _2241_ VPWR VGND sg13g2_inv_4
X_4626_ _1575_ _1327_ _1237_ _1313_ _1238_ VPWR VGND sg13g2_a22oi_1
Xhold510 ppwm_i.u_ppwm.u_ex.cmp_flag_q VPWR VGND net1162 sg13g2_dlygate4sd3_1
Xhold543 _0090_ VPWR VGND net1195 sg13g2_dlygate4sd3_1
Xhold532 ppwm_i.u_ppwm.global_counter\[6\] VPWR VGND net1184 sg13g2_dlygate4sd3_1
X_4557_ _1225_ _1506_ _1507_ VPWR VGND sg13g2_and2_1
Xhold521 ppwm_i.u_ppwm.u_ex.reg_value_q\[0\] VPWR VGND net1173 sg13g2_dlygate4sd3_1
XFILLER_1_229 VPWR VGND sg13g2_fill_2
X_4488_ _1329_ _1333_ _1439_ VPWR VGND _1289_ sg13g2_nand3b_1
X_3508_ VGND VPWR ppwm_i.u_ppwm.global_counter\[12\] net594 _0682_ _0681_ sg13g2_a21oi_1
XFILLER_44_1021 VPWR VGND sg13g2_decap_8
X_3439_ _0613_ _0611_ _2255_ _0615_ VPWR VGND sg13g2_a21o_1
X_5109_ _2047_ _2048_ _2049_ VPWR VGND sg13g2_and2_1
XFILLER_26_642 VPWR VGND sg13g2_fill_1
XFILLER_41_634 VPWR VGND sg13g2_fill_1
XFILLER_13_303 VPWR VGND sg13g2_fill_1
XFILLER_13_325 VPWR VGND sg13g2_fill_1
XFILLER_14_859 VPWR VGND sg13g2_decap_8
XFILLER_41_689 VPWR VGND sg13g2_decap_8
XFILLER_40_166 VPWR VGND sg13g2_decap_8
XFILLER_5_513 VPWR VGND sg13g2_decap_8
XFILLER_5_502 VPWR VGND sg13g2_decap_4
Xoutput6 net6 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_48_255 VPWR VGND sg13g2_decap_4
X_5497__281 VPWR VGND net281 sg13g2_tiehi
XFILLER_17_675 VPWR VGND sg13g2_decap_8
XFILLER_32_645 VPWR VGND sg13g2_fill_1
XFILLER_20_818 VPWR VGND sg13g2_decap_8
X_3790_ VGND VPWR _2224_ net661 _0114_ _0923_ sg13g2_a21oi_1
X_2810_ VPWR _2164_ net500 VGND sg13g2_inv_1
XFILLER_9_874 VPWR VGND sg13g2_decap_8
X_5460_ net46 VGND VPWR net936 ppwm_i.u_ppwm.u_mem.programming clknet_leaf_11_clk
+ sg13g2_dfrbpq_2
XFILLER_8_395 VPWR VGND sg13g2_fill_2
XFILLER_8_384 VPWR VGND sg13g2_fill_1
X_4411_ _1288_ _1298_ _1363_ VPWR VGND sg13g2_nor2_2
X_5391_ net270 VGND VPWR net408 ppwm_i.u_ppwm.u_mem.memory\[50\] clknet_leaf_24_clk
+ sg13g2_dfrbpq_1
X_4342_ _1292_ _1293_ _1295_ VPWR VGND sg13g2_nor2_2
X_4273_ net739 net764 _1226_ VPWR VGND sg13g2_nor2_2
XFILLER_39_200 VPWR VGND sg13g2_fill_1
X_3224_ _0426_ net812 _0425_ VPWR VGND sg13g2_nand2_1
.ends

